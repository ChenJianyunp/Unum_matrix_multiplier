`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RKvPotahVX0W0xVgAVPpEpW3UazKOPqmIFUllrqt+iSZHYZgtjk8yNjZieS2izfS43AOfK6rW58p
vX9zoz7Y6vcqKYAg7wn4zKRpmYB8qij9KIDIx5hf5eFitV9Up2xWQrGhAt/CJ+q2h3srIbDboqoA
5c6O0d9RYMNRwFQJkcCmVBi1wYyz/OXFpyMuktnsjgKBSQNuYpO+/dizxap5zs+1orCFHIi+DM6Q
r2NGFunfCGP8orCurg+EXnokrK3BRpHgJonBMZ/4aMuxHpzB4z/bJ8JZARgLaAd0duP3f4R60nY9
df3tmlAobSVLHYPQDL+WgNJIAjOmH4iDgNSr5Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19920)
`protect data_block
NzwTZfbeqsVdg5St+xLO+2dCHI2cO4987rA5W4bezIrOoloeqU5Nq9VNISa6mnkEVTdOQsw/jHFX
rU6PTkDdHjHPUB1scaly8aqppNYrYWJnaJA9tWnN22ruDEk2Eo5EuIQYStRylB1sw5jhd3XzAns0
hKlOSweVU81fFyeVsGUNf5Rx6VX+QtA8Vj/VMS6UdVF1/PH31L5N0aGDzEND81A9dDeLA/DMMFbs
jKVf2v1KYwW9AQvhf4As0kiDOr0vtqhrKzu9mOyCafBGzq9HNdicNdSYpDxUg1NczuIXtAVvLspJ
uKB4XJhX4KnnQpPYZSQVz12aNaHaHuZMBS/Lph3mSQfk+QN6E7jQatYoacLKBm8FUz1qcuXPIH2S
+5HFIsRJaFYZsNyi5EGf2Z9GcWE07WsO+nsX+Nxzx5cwxATA9m1tuT2aOSm7P9Z3DEmqAQdBMgCc
twPEEOXU+ZQmYUeVlT79ZPijmcnwI7mHCxx1dZsaNgyL0+849z761GR03FaEaa1H7zT9IziruLp+
4jLaMkfBhwEMrI8pUVKJsKCq9gMFKLWXKNxTg1iHtYoO1WlntsSl1Uk5v32yf2Oxl8cy0NXNMnHe
CMb4jSOrMk/TRmcsTcPM1sao0wvfZEtb0G+9MDdhFBbViRErNgaNdUjSlxReWBISV2Al0dLedxF9
c6rDlRlAwMyVRr8/x+ryxHRYT7QK2GMvjMgL6XNB7RG/YFFfHFsg0yif44gFjm1j3F7muwu6YMEv
fmkywY1G3fqDakBIH8lejn3eEMgue6CY1/K4F+dXbsF5xwmmcujxSwQZMI80ichV0TfH1DPxkEUn
wwdVoEpmL/TMNIRDGlIeAjXKePAHQIjdtCLl6Jox9CGOJggl7D8yKKDMmEZ4dT/kMgEtRVMb82kd
LPBRnqyu1pV4NoI3KraOVfsiVeFOs3n2iAlp7fIPcyYYSsbpxRJMN8O6pmOlbfITpfZIu2/qIPhq
xHlu4gXL0pBtYpyWL7snpp51rgM96N6q29iPK5D6YfnVgyA8pQjYtyPX+JtkWBr3zOwKkm5gEwg7
fad8ZeVKUaGLzWY7fl0fGxzJfvVNJS4QuVdQ95LfTSZCi0+iZ+0gvXiqHaQ6Yrkl8mSyjhfZhRhw
mEU39KAtWMawPuWWO75cbe5Gy4qcgkW+G/xxGbwzLeRKYr/mhzMg0JMaIBs585q/9v6yr2b+Hv7D
/BZ51vNGb6B+guQVELLXU7qo8zAu+M85et793k9wkoONX89vTK0lzHX6nt3RvIEHwGqUTRQBdaxY
pP/peyic654wSrUqDZHnGkUEBuNz7xDTt3zJ+qrpBXcHmAw+8bKsoxiOslPQI6Hw1H/ZUBwhGKKP
2t1ppEPBHlR/B5pAgOSpw03Wvo2No7kXGQHvoP1Q2soYCb+zwlFQqQQrHXJtdK4QcHzmLeb5jOMP
y5XxfnJ/gCguopR7+PGGCeE2RNJKYu2OuO+oeiR1EefhHT6dSI3/dzUi75Cm4PzmS0vr6lOoGuLi
GpHhwd4VwMQ5ZyaNLjnivOWTNPti4Fz5GQIACXb6blRLeFGmh3/uCE1e5UzeHaW+g635UPn0t/5b
WEAyFBuBi69uker9X5DPjtJvzn/UH6Lx0YlJHvcVsTACuk2mAJPPb3r3GShBpuJmZ+tSSnpvKB1e
AvU6qqHUVqJRi8M7tqdbN1y7CiIXSKKw9sQFXOC2EowlgNNMzowLfN5XudwjUHCMSX9eb77baa8B
EHGHZttDQPfDBc6LJ0QoCGNhmxljkVdu1r6BHs53u+nZYTPXBR+kbPIAZRcRpGTPnwFU61+3SSQR
KmQvGADrZ/Um3nCFvID+VFKkip85oesamhNxQmApJoTGuwVC+uW3jumpUlp2YsNtntiI/WfLUsey
CyctfMJbfjPBVawi9gsHqRWp61pXURmRJKn6Sk84g8NzJvZExTcJUZt0kkaLovmM11JPo3yOCOCI
ji7FCI/qZ6E+R5raFmor0HlnTgQznOK5ttM9YjyAnKKyrFWf4pQg3AxlicDwBXuT62MH7GPXX6Ml
aeLq4ctjgeOTtkwKAI+087XXLtukvng+pkO2pPliCOAcYLQqCukW0Q9WJvMvYmSs9Zd7ii/FQzQh
9/bk0D7IFXizHXOdTXJhWl9cMJb5VDbT7pfs2xYmgd+ggWrUWhpTQAsrCxfG3F/lEa7XWIpQN//s
uyqqgCh2uLDZJjssXO77DsOv7zKaMqi5RzqYXgbYxIMJJlHY37xFV0rwrtKOoalc5NaW2FOnv86J
P7kx540A++ts9unOYv8WMFnPoedX318f0lWlygJNzJv6PUo2fxQ6EV5d7kRLD7NHz6mmnTwRFr3G
mC5ZIBtYImF+8yUsn2Gy0r6xb8m86R3yzmt1Du95pyw3ZmYwj77tmNIga78aIQG/26C7zjl2OM0B
YM1M0aEAjnrOy2F8jyHLG2jNJYOgA3eq8Qaf4KAioj/Bgz7wKntZK7XeAH+911asg950nk2MIRor
yiZWH/6KgRQK82pIHR+HhEfKexbQK0RBicXXYizFF/Tv9xxvWsFTou9SpkutVgwZDd7muF0tGGbK
HfH24TX9I1J2N0ZWHb+A7Owo4DxGi7yjL3yJlauGM+P95aGUBBWoDF+amlt6QBc+Vl9ECmh4umru
2mSYUhEnJ6fJEWprzDt23UnI5Yaqni5RkIpb1kqvNUgT035+174BtDcCTvnCu84Foqy+q8iTDlTH
VvjUCJMKiDf3GYkX8d7KHRsoXaZZVWkLUKS/MG9KJ9xDgjm0m0CtlFYd62Ptz9o/5Ev7xDojU77j
pvVvEuTjkoT3IZumAIVFUaMkEXpQD0Pti/+nxNJ2+zVy+fImR0KbKiELE/T5KoJwZUj3BccAOtwD
pHcZrEjB+GAyFw5QGQgxGYUTtkpqC6xwG4hq5zafIisGRCSyfg4fsduSj426w7v4mmkFQ72OTBqQ
hkaE+pqLypgDEO/f33sz4Z5/eISYWOqKZPpiw/eY4yFQCDk6UmyGzQJIoOsp1YwvvQ7q2OLakOmC
NTI6h5NN9I/Ng0pt/uzM4ZcT8+rA3VuHKsCfciztf3YZB7w4n+nhKoifDQmK+NVqmPREkkNg3A9t
KBXDwmDqvgqn4mrc2gZDwcgmrhV3sburmh7iOVBeenK6rKF6HsfeOBBBIRWLOVUFG8a2VIc3sOm+
4zGjMWqrCH53Zpf8MjT98UV2i9Sqi+vG5tpj3a0Bu4xtbW8/Gb0J9fxAURVwLGPTPyYnsIgCgGb7
PJyJB6kVLfbm7ICa6vU/UiZcuwDdTnqYyQSHvMKR4Pppt2XcNIeYGz6ubQba27/gs535Me5CJy5o
rNTpRuz1i8EYb3l7LPFYtMR2GdWFyBqd6Or5F4LQM5JsouWvuTIzmAUxdRzdom1C5OkPwkfiK3fk
hslZTAw1g0bzb38vwc7aCxv1Q2QzlhC/MGWXZ6N2Yb87sfZbRctbDqBta09a3olB3DlZldd31Qjf
lfMCJGxSkEkD0g+CjitmvPhekQCrToKO+qJW8tKiiL/nNKSJYsDKG5lSGlFBCtEF+PyrVLufBMvO
bqSjMOMIP8EsOYKFs5y0PDNSPTffK0L5q09megLnb4a6IRa0GjcdOa1yZ5JX3oz/L70mlbXMLbRe
uUq0BW9i6YXPXQK+aEVmElKbCbFMYnIEW19lIpFMaaLOQRMFHh1tCrKjSxT9ocX3dPxxZfBXtXhN
tK660C/TxfPBH09XJYG3AmH1I6hOYICNMZ36LVmTtPb1nhJjsF5ixEzyCfnB2HsdP2ZyQTNuODAQ
E5xBhTNfdoG1pCh9Mpw0jCHzxeTSoDWDX9ou8PI6btBZDrsq8sG83/fXka2V1M6hTiYSHh01vJ90
nsmj8V/+aFe/tM4vEPvRb5xuJRVTkoGWWUxPewbLTu2JvgNpFfAeYfJTcHUYxz3g1sK7mkTKTuyH
rtvJzwcH8r3kUtiwqq8UfciPDQHFlA1Fzno+BZzPUWEPx3XuHz5YjAf53QkxZhlpJZjHrlRcWTZ7
KMVTeqIvB196oT4jXBGASx7z76Xgq6uibBL2Cc7/aVj/+1rzsS4vLeyk7xAYtlQn/xWX1+hGL85L
TLWb17o9sOr7XT/4xht89cec7nLC5FuVEeOP7cX7gR2daffE/FVDhQUwtLr4z6652YfAAb6VtpZZ
hv7fm22w871X+Q6K/5rzBeKk0qowwb6l/cUD4BAwnqHSmCi8i0vdVFtL5+VlKecZHhtxOgI2YYsi
BINgkYOwQj/J507lr7SpREgkwdpYuuOrErHb1nAkYe46QbMffmDDewO5WBRdUBZ6gBNgpIrGULqF
WJ+MjsfdJ6n9ZIAVNZ94mvhW6kFPTgkjyAxbwXv98sWOVsR09ix651Dcz+Dtnn11ijUqZTBZb5kD
JGD95vSJDAKnTf7Vw5M1XQOjC8/v2/Ha8IoOIm/ojHrvznLBoQRyhzC6XByKfAsKtg0BE/0uUEpS
XXMw56NB8V2qgQu8XDsVapnk9cElI0ZwkN4bBbPLfuAelTzBry/3l4P7tKRVBz++isiSrdx+OL87
UyNr40f+e+NelV4dwnO3wM8ekPZbtA3t+4wc9eEAlB0jWN3sY5NMV6VsADR3flIXIHM6kjkfyJG7
TY09qiOFUhCjm6wXyTIYMMTrNocWbK3l2CJIooV+yHLULzbXoxM2c8JT01B38BRMc6Sfnfo3CCQB
NklpMypV+o0S+K7UfW6k3b0uAUmSSOZEk/8X+r0qSYONMqkL+9LrWhnMULRLx4V+LV4O4xzFyfMo
vIVmOTBP0SpZ5lK0dQbmGJGT0at6LYzYxG9EAaJdv2HsKwLkIBGFxAalsARZjdTYSThc6wiAwadG
IHzpCqUZDYLgrp8mvQRq1Xx5iny6hX3sIxBZaGpwH0iVo0wTaSXdYOyKS99XkVMMsbkAsNP120mS
75VXj3SuD20gLgaYRlvkacZyiYAhjIR6fK6Kt03XKsEY1mAWonGhLS9qv/CVoWTFKAWiBYBuHU5W
1fw3OX7PoHOW+WcJn8Qpqk/JAG69IHjJsIl4aIyvKGTajHYWGcU35QgDkxxwXOFzdiH10W/pi91l
wfsuvmfbyZN+XAjpjRMvzT9Cy6jwlrJDvXBvJHIsRu04i1DKZnbInLoPcxX7FM2N0P/HRTuHLWA7
dhRAuqvFADQxglgaa1dL7q6SsRfpXfk+FJ2qir+wJBJwTE+H54eJSyKOqsa+Q//wyjixBC2emhpV
Mqi5wZGAuS5UxMLf9Gm/loAUc5Z5aBtz90/w1ohe07qBDNufihWLnt//v4RyKL5E60C+/7wA02NU
02WB5BV9ie6A5ygQqDG5bjX8LkBHRuN5tRoWUZqqYit6X+mWVyX+DnVlnJkcg9qbDMiZqI9tHzUQ
ECwlV4BK9sfwLtsCwd6Zk/usIEEprVPJJ+OvriglQBTS2EaK7uqYy0OVjxrlEZ88WCfWILYgkbDV
z86k9Evv8Hhb4DqptnpnMIXe/haSzqtWY/HuOyBCnXaU0uIXk8QdT+/VS/YX+TV3xl0gTWEOcnkx
gShm3VzlssyLKY8CM+/ay8pgc4gdUFZfnyo9QzRMwXkW+Q+mzpp0OgqZwz9fNNChISYa9yz5q4NQ
UCPOHYkVXBv5rfZPN4RM6CSz4qyvmWt6+voeWiM1B+Q4KJI9tH8bSTuTiKIRGS8HbNZjkXJVcG/h
OjCXhNBLcG1gBrxvK+1EZ0Gl5v8kJ009kTpBsBrB1rCub6VYdHT1KglQzZELZR17fCGjJRvp5UMU
kuEQkuLDQau/42qiq6UfYDz/uxDSt8d0CRXG3Mk+/GD7plB62smQo08yo1OnwrNhVtbukUf542Gx
g5b5k9fJEIWDh4DEMRTZxzdt5fE9z8f9MItfYmHFdtlVqyLXKhPUWboWKPyybT+vvLXgn+HmZxP7
LShIfHRj9wAtzu+0fte82OV2B2acrDGyAfeVghxwQNx+HcAEHCq2QLqPZTkoSGevoLg/dU6jpWzi
9tXbKSfNIHyjGCYeAWhP4alcwlZD3bsnSxaAWZLEg8fAzDst8n05eazVX4f1Of3q18WOpnZ4XJOX
FSEaQQ5GSthP/rkXkocPLtePsw0csWTxaCWrBAGm35CYiI9+0bKHaIJaj8lcygHxbknhcM16v0wF
7Q9iF4jE2zBEKY/4u4Y81orYEcUInbH9PPHYG1h0ebzUbxwLHboc2UC5xqpfYYMrlpTbtzQoqSxl
nsFWGWwQ+nguZ8V2f5VxBVoxPl6+uNriGwiOhOHigmMUy8IcH//apzLfJbXmvqH2sgN636CH6Ylu
L/YJy+eb6kpwWPdry+WOyZT0MWtcd1H+cZ+hEUivLIyL5/6ccBuNA/KoqK3ppHwSO0Ld7T2BmXFz
RpMKd562hF0SiXSHTW5XUjztLpXnWBqscpZptfhmuGS1EiN3uIUCd87D3Ti8TtUo3VJFxQxLkFxl
Mh4bOlE8ZqgAd79A635WgeoNozKUoN9ppRA7JwdYEoL0zk4xbEag94ymRBnv1Ysy3PrLHn+bt+KA
SdjvmefJQh+T3dIXGOYbb15rg8DtVWsaDq7UBCrQthQl+VzRWwGVWUU+N0K5H9dUYgsQnWyKX2fD
khZN3jfvubiBoYfgCLBRyaamE0qQfp6IooRJ6enH8znNJoa+kUjqVkB9wC2tvAy6YQVgoXJi+9Gb
A7fJ/BFyxdIoOEZ0JHZe1Xd8/9feCitpmB9HwvwaV6mGkAKLoZdQTNFN5Jclo99Vgr04oQTrQ8lw
Btoz3YoR6gJG1DVM9ND0rT6MCRHd0Pi1TsozaTu14XdRvxX+zOOCrF++wPtAI+GIgri1UXSprMmg
fPOZG11cQvUCKmE+oHltmbLWovHOMBqF7ZRkrH+RwN8v/uKT94SlnsEJP8nDHYZKuB5+dN+ZAptu
We1VuvpFyuyN3LRpLim6xB+yzYi2XtLALJ2FiNKEdJUC7a/GxozatLJHE/QfhiQMbMtdKXP/TGu3
HnJGn12cEh4HMzDvN4SnADdh6Gga5zqnxV/Ak5ykdyqCcdC536yn90ID1+1ftuDh2p2VRrewVjAW
Q6TB57uKSLAXuHYXVZ45StA4xbSQDxZy70j+UY3nN920LwuJpek35JFBund4wSV0bRzsBDJMR+u1
l57VP8DKgh66wO6p0ucyKtuJU2Lb/j7bJkFfaEJe61rJE2pbHXJC2vFxPYZl+FtqNb1Z3xAebf8I
rhPPQ+lpw1nl2N1SYn3crXXU5JalgIho/FiQ2equhj3mN02IRdJdp0HyTfGjXM+RRCAB0VngMO4e
B/ksQYpUT492ksr8iAMmZCoHwk90qJR/JIQ5SauSH1iAHBFUDeEIbKUFbh7c5ZsVydXIsGMwTdBD
dfGfMDSBY7e51IN23MRAb75jF7fnzHat0zU8wP7VtVsOyof1Tjza1KA6VOk6sIc2jvH+jYxcwztf
WfVrB8xvPEW34I0487I62b8w870ZWIn93oongrlgJaV0S3ro+C1igjPrXHKGrZDGap/6dKjiYuYd
8LxspSCpwxFD3DMV48/ugwXX1LoWl9VCU8ptAJ6B2aUBLIKwG0Wi3oXHmYdNUSyxViubc0RqjcIj
WpptOu7qEPixag9x7KdgOGz2o7WuwoD1R1q202d8o+jbIC3NQW/TmRmpdUFsRHEdQne8vL5T1JGZ
XB/3M9JVxub3eDOQtMEqlCR0x7yVAMvrsH+7gq50lqlkd/tNVDJa4KfGTRtCA8gCAEfxzsNVu6cf
Rg0mFgASdYYKY1AV0SGZy+faetLYvx60NJadDvGrvYdwtB7yrzmAensM8OSgmn1a6/02yi6eNYd7
cRIHzkGO9KrtjhELVtHmqN0AwVFKXV9/KD7ZC8T3sensOj/zZtjDaryIWfWs0J+l7T8MG8Et+ri7
JOBBh5OhsohCT0GXPJohUuSta/9c/Z45KPpyuDdLcYG1ebut6XacMY2AOhmTXkQZNt8Q6G0evKTy
mM2MVC/yDNnK0Ea4GpLNyv3aZo8DB0nY8MwHvKU0/7ozDFP/jbJ1EJs1Hbc7o21YUU7/f6yveAlG
GEhfNL+e4hRgu3mNQ3XN41/DGv/AUE7OMgj5j0oXPuk5whVlZD7hMCqOISK99ou2DtwtoDm5Ylpl
MNCIzoZaZFXbFFZ7EVotDImpsE+noKU8e65t7EsJH4sUzBUD/DDaQu8+kYFJ2VP3HI0dcTqX9RRz
PxG+yOXkvCAIuXc5SDUOnQq+W/+CwP9qpL3NiNbhDzc6YyJBRdLLMVXmPLekTqkKVYbZNLXnP0bS
NMiLrR2PoPiH/Lk9dghiG2dY8Fg4obmDAH8DlIgLL2wZtEjT/XYsuMoHjBEosTKQ993d3bEUkEVz
lI547T9H97CeXMEiRc2kF5EFTAW+4p+qoFAjSqPsXkqjqkYL95eZWBBESaossQRg865BHNRYP8vP
4E7XLxPwAbwyh9ME/L5MPE8apRS68tUa+71Ug665QwAbJ+1DOeIM2378ALNdDiq9++fKntxwC/IX
z6MDUot3AcPu7OK4XMWphcZCqQOR7d5BbEPYpTacxcc5pH6vxZY78hMzBDVWaeBrx8Q6RrKzGShS
/6DMa674UzYYfxaJtu/f9XSz39q/1ZsD6Bm/uPNo6dqgPUC626KELMJUoHLQC51qpytRREGDoUeo
nrzYXc3XjDeraVxieGN1nZAfaZsy0y/cNS6pUk3MIdObdQl7R+GoyLBEwc/s8WkuHOG/A+qsiwvn
vfTmYFfjwYLDxDDmOe7SPAClL9ExBqWRvI6P0JwcK4rpW4K9PL9RYI6k88MNRbIcZEuJVSNNaTMN
syYppwgf9SM6A/DfNUYiuHEI7TpLkDBhLZ7IsXeqtgZcw54RooLBZzmyF3z0cOwctyF3UMoTV/XV
jKn+w/4Ehv/CNbwr2y1lT30e+osjCIS9B3JPXi5UOShlr86CQYSkCNgxb5+gaNgemKbZWyM8/yjD
yJHcMrIg5mHpt80EwsDRL2vYW2ZdVsLvUWU5TGI61e87Q9slOHolrq4tiiwBFpPzLL56vDeMQnO2
pBnYcz9LIfwe+TjANfmHxW81dkHYilkE0YYaWkfsK8rjCwKjx3+oFD9tyUSqkSLwhRd5pMpugHrn
K3kQ8yudY0KVyi7mfem+TLY7xH3gwgaHrv3rSFraAM/O38/1URtAHUf2IEGxpiNxOjS6PvdLBuNd
DwiwVycFZZ9XcQ+jRVVrJ3bbOwnDZEC9lCGBB13IpMLBnHBjJa1s4eLiRTF1G7IFKP8njH6VSXZc
qqJZ6n/4INbmvldZyvkffq9Fi3NTOgzHlmgZAdmyGc6C70oonoFu3OHu6GPRfOhuRDLp1V8Rg2M2
oX/gGKE0bLxdBg2rDbdO71C83CIYJsMu7idoZCq5sFwLatKey9kKRIJCdTdQStFQEY7+CQiLd9pK
IC4tIaNxJorYN3xh7Hf4N7PpYxeSTnKhzGaqZLnck9NJy9ezMCgy4AlUq4sRWBTVrj66Xu3BHRzx
Y2Evr0HlC0fNSbRots8x/WcSdX8iMNckTji5XvqdTCCiDdrIgg/Uhh9yMETD27aNFHr/+m1FY8pU
6nYh0M39UR+w1YeVghleXAIdVTfxKSta300JpnSAjzX85vFPD6ODMy1DdKXyMd+PkALyb89fKNek
L/qdNLybbMVcYAzleoHLTADJ/zHbe3Loi5MqMD31mJznlRjH3V8Z2dt6YAsBKMUlPFxo+SN/m05z
9P1SpCQVhMIl8o3UPQItcyiEJDsG4LACl3DZeQXJvQXIPhJrf26zWHacxKum710CSiL/+HOCMjVt
ja81HQ5fKs3NNtKS6wJNIHQXxMAwgiIK3PfKX8Ej/ZGMiv6UXbYmsquQwezMRmjIIoduu68L7FwY
Rp8KFA7S9JHAdAPtRi/1aH14uYpclP18yfizG3r2RWbv5QnxXktvH9ttw2ylIIqXAvD3pxDtXAdL
IesUp7eyVhWSxKLJcN1REbJGfTF/sSvYPcjfiypwi6zE8W9J2QMgCTrVCcMtwXSvt+uQAeynlDAb
14MEZlxFtT/j9HhZVG9neojM5815kgyKkLBuf4GnABjQoru5WYwkm3TFSUuHoJO6j/YzrpzNCF6X
w6gkF1GxfRzqp9A8VNWxER6Uex9kYwEL3TL1tcXcKXajMpd5+RbPI+xpvcEe24Ibe/YynlOvwSuH
lSNcdxzstFusrIUclMqHScun1PXQo2dCbsQFXQ6ul+fHKm8IEvRcqJLG6ZxCIO2J/tSBSFkD0cWI
ncUbCQhoD4snoUSwzuVGmhnvCTb8zlxr3X8KJPhVjJahmhlEv8sEa6aq4rda7z5Z5rsMtEPeew15
zQXDmwZMp5QlZHCas9p1tF+2V8QUiavRcstbOKuwuffuh2krfneFkzxbljw6ztYMamflHAsgHMxJ
0HZRPmCHqjhOJfcMxgXLwWLrBbcbwnpr/tDNDf4h5GUhKfv7TgM+RQooFu7DsNOd1sjAUja6WUEC
OQ0cU6NZ0rF7DNnG3MNneJFacq4QvOePfFpX0Ew9ZWmMDpTcfKvG1L5/F5pSofQp3nIBpRxJkwt7
/WorfEwnwMevQG4hIlpyuvGVSLfsN+wQ5BR5llU0NGFm66mTnt239e+phCDeU+EzXKhlLjzr/Cj+
W3nRfrC9Dk/XWKqvd0oO2HOk904JOy1/nrXNogNgsnnMq8a/3PjJ00XVWD5V9zqaFErII/fBQWfd
iCHZ5ERv2+mRp3TU3FOp8Ig9n+couA3o6Ko+EI03rzeya4X3IBSpADG2gwddC1/5XUXMpYwAlOaN
HksRsPm3HvQ2vY8C1X+cLNWm19vxEwUscXIiBXas/RPwKwvWQudD+Uq7aK287MdbykHW/84NlCND
iNz5HGtudn+rMplBwXV2MrVA/cdel/A8xHz6o+I9Pne5GkF4aESPVOIPpTfFaiQd7hmLseNn0qk9
sPNrEQQ/nap8dJ+ufZayD0aWKJIiSbXKm+F0bkKPVOmKdbzfg7HYhQ0W4sl8QEtNAXHdW3/Hi/vO
whk5X87MbWU4e0qd48gLsIpYLFq2Mr7wlAlDSR9560H2eXeeCyHyZXqZoWxf0gRoe640IvL2Yrwu
jYXUIIa9iqAW/2K4VHHYTisgLhxSva9Jc9GtSYHOUJK9nWVjqk35204CetubDWqimCKfdto0733s
z1VsP7WvLlp2RhcZ0AXdaFV3bs9bmHPgdJwKn8p/L/SjpyhxZevdstIiAr9a3r+dFKwD0qN3PT45
19q3lOTk3AVDDJu+0MQPak5YfQ9OKXOwEpxy8WV+FtPzi9yzWZBzqMExpaAapHJc84rUobmD2tiZ
dwk00oUU8WI3O3RE6oTQClL36674PtJimKuKPtQM0TVyLGjnTsOja4LANeoJYSeOw/veuQkDyUP0
ahdb3SOCEg1zQy6oPNJ1kIE1eYNRttNpD9vY/a0UdKjgx540WgDXT4F8jqeuQKaw3Lapjgk2oxU2
vXF+IWdiaj1ff+IhYzbnwShbC/ECwylJv06EVEd7SdtT67+uG1aD7yMcMIyZF9srA581X9FFzKGa
pKwGjjoG5KV2kob/F5Lhgs/0jYqte8jZdnbam339sYtzrhlK1puE3CmpdOMobcx9j8qRoJY5+4Jp
CGaBGgWe0cTDvnD5srMTGUL4R95VaTr5qV/OQE2BkjMsQXf7m049mT98Nut/dnX2mmCefjF9yQGN
Le54FASAM32wTaTjjVzzOwlLC/ogmmKZI6e576OigmnQr/19SYukSeFj+i5o/JBoNFf3OXvtfjzx
vvcQyyIIqyK/TTo27X2Qu4haaX3U1qWdgKwlOO2WnbFX4K7szKxa4hj1X8IXn/snmXr3tF8AbPIc
nvDwOCUys+YUStEBK04VmxkaYXBRDYTtIp7DoHxYIVwEY2Vjo1ItcBXDXSIDS22FdUIwBCB5vPBw
UuHW+0ZXPw4WXPCOcXlLer1lexhZOmkgIJKwZw/mr3b9IXARAQu0+EKiWE5R0vy7wq0ngohVjJ54
7IM/5/TE3vSnun8Jk9ygJZEKY6IBEqLq9Ybe1muvuHSSyG0sj2e4w0NoeaMnE8DhRspGiV8pgMxA
sOY4EFB2ApugRBuEFgNHj+/H5bK35FGB/3poTfROEU/Q84wqmWAEtDm/1W9XKM+n01+lpqFQ71qU
4terZ3hso+OAyofq6uCUOxHd6G5HVp/OcJKhAB44tWXnyp8X9Lp+/w0pHNt1VikRsG8nHU3ydLwR
3i+NbHYhpH0Sk3kWLlTBvmrJfvCiFvcxaL8JaoR573unqVIqdlTxw7kzN5QXl1o6rG+o1ACPl6jy
+gFZ27ncazpG1qzOyzGWXqDx46MKbxXNZFFjSKN1y20ajVYWxRozA0e9o9ctujjLGFjoOwa8eZaC
RzVjmeVueCBh4xpuBzMHAr00m5GPYyT1997wdfiawMK2SZWwBeCqikHmNmp1dik3MuBgzlJvH5po
Jy9HdE/xtH5ShIYVNFF3QNqCm2JC14Zp1hhocsp2UfuagUb6iReYdl8kBFUSBF04fy/dMXdN8atc
BZaGZhx3vVnAAph8qWNs+d17ESB0EOBEZ7BfVDrZVretMk4sVvSX2nHkD8QX4TpnXK0+XrvAAkNd
SDwYvFCLanxmSDzZv25tNfw6lxCcC4/rxNeUl1tLhZlw6vHufWoEbVaEzABE37SmuXQw8kQ0uYx0
6x0ao/6imx/WKFbtfGAP5Yz1KillCScYHoUG/3XchYTDEHwgtt1ZhWbKbTXVwT3nhw+VLoU+/U/7
jjpzGeAdF/n9mV16ryPkP6SSZ6uNJhLgVl7DJYi3HbdGgy40axqEY1+biJAAtMm3woCHsAPDYMBY
Id9KKke9r5O1OY1mVwFB5cz5ZcDiL0BusGcNfZy6C9b/xKN8j0jEoDQlpP/QRpXIHynQW+PUqRxh
ixdntjX34TAFNcjI0wmUjgORmDzSYTYBPkpWz0g9GazoDzjdA4afbeu/pld5ycAT4pbqyqOCQAuM
k/PcbM8XHQK2bZbcQT7yaNMGI7kMNxfiUfyXBpp9YA5CLXL5yeL8T8V9ORgOLh1R0PQOwmpHtfKz
+iZ0g4V/L1BH1BUsri+8fCvNiT5MNFoDVuinyIUf17fq5gZe/8iqnzvopyWGuIR2LUUFe3ImI3c+
ipYumf05OVasszfPrXZ+T3+6cfiUMjY2i6O7Z3zisqyC6w4K29gLmcA+J4mlI++Wd6X0dRYpnOTZ
TuUoIxfqN7lVNMFvgBSlmjtHO+wpLPhY+hcpEaK4M1sIZCUUSeoo94t5OePF4dbm/65RjBbhT5Pz
1DgZcIYAzKZXbWjdA0dZcGIyXKWQi4F0lJ/q28YMtSdbfku/udNh7OCT6dkLUjSdrS+s5052EITB
joClDpbAuBJLl3DQfpMuSX49/YcfKbyt1Brl99w3gOUfVhp5GwnsRjrFtKhp2pwJ93+SjnkvxsED
hej/uwp/t90x9rDecX2I161NLjKNArDNYTBJmnePNOHHqdKdble7dA0jRo6Vjv1u4Pza9/CekDHX
STpDf/QjxBae5G/LLlxkBtyRC/3NJvpkU73ODQx6UAEGnhWwS2R4iDpnIbjxR6l3oZ/k26/m9jVs
Qa+CDjtfTtDUXkwz+mv0xIYE30Qz4RAeScwkuQNCaA/h72LAkAxBBxuFT5NrLDy8gRciJ7Ox+KlX
V3/qlBu77kzSAmGEgTD0FChBUyBFfRtYBQjMnoIXl6h25Gjn/2E5LG2SRO5tGPxxbIy5r+mbnklw
vG2/Eo63dVjpBGZjtlpxQ5E/1DTvoYGvXDmaavZyrkpQa0PfjGdyAe6n+aV8PdfydB0uofmvYECQ
ips8auL6RkKQEu54mE8IiHhOyW8hbvSkhr5zOIvOmZwDuvibTx9uDSYuNFMhuy1FySAlU4Mxv+gq
UihqGuxoZzw5iWFadzH67pTKT8rQLznSDsh0i/CW27QbaVR6YSJOYHLIOvPa7BBc5OLx76/1uHHd
OBzI1CVT1EP690ikEt2bn9/ZlTRxZ5X3q+u1mPcr+iVaUPAVPy5qv0YTvwbhISnzTE22O9WdcXDm
bPDwDFk/o83YNJkGQREDXlgPLd05578VAd1zSt26yNeduwkpgyq+asKJKacR24QplY5F856/P+2O
pFK3E4vKzxIbOfJwcnqkT9yv0IcPJX9oYVFETEhKf+2o0c6gr5thI75f/RuiPqOqIavBGY/9WiDv
hhCaauXUzWC8REgJbB6a5nhCYo9hnw6KP5YPfd6Zde+Ad1rmzt01Cx0LRxXoWO0hHhiV7iPQGh+6
LYGEjKMAIGH1S5JShAnMCHII9u2Cgo5qNNW6ONd/qGsf0MC8OsfHv89CT4uLR9eIqy/SOLK6wcm+
xQfPrGRf3+7rnzuZeE0io3UgsEVR3jX+q+Y0uhnKKx0bLeuIgki2bxbIar39fshPOJhfwE/FWDYd
6kJiXkrueN7i/TYj4hacm4Di/Rp68ObanbUqf6Nsv9ihY+zFYxUf0M2VGKInSgdri+UGxqRTjdCO
2f6qFGiFIkxHXZafdZgcuWRrynAXCE12mE7p4AomdjGMKWAHwdJklez7L6Y7S0dvv6LltQ7hZZr3
m861CRGR1V+jL57FqoKgSI++2xgguZT3QwGDppdGnihqDkEmIGtgz83vIHFY8UaOlfMtFwBUHY1O
ydDKv2yMI2trtMtasM3BsW4bGoJTuGIlfvO+YOjKdUKBQXg6m1k8tYVQJ1t12U0TvR2NrU6O1aq3
xtgnKpMKYs8SOG7vDfrs4RS0UDQh3a/X/qX+YNDfq9IsdtMP6gf1XkObuaswyNZOT32UNYq68IeZ
IuIMX8f2FcXGfkNFnHt7B2fkehfLGu2PFst1cq+fP9J/I3SzoH1QCm6817WoGf65QEdMu5FdpTFl
dFRKJ59CqRCh5C+9RRwyZOKYpIlpVI51hZDSKUktpm9fmy/OM3Xkmhl5TdXF/93o9AaCsuqaNpDj
7DgXjwydbNRr/aeA4HZn8qVDj9HW5aXmHWHtvDt2lqbOUrvJRCs6HwSoNrL2asH40LOgCYyqna8q
avN/yXRvefDqGp9cVLF9XdRxweaJzP1q5WXao53cDC3FAm0fBPu3sugYav1B4j+Yf/dKz2XJiqkm
QRCMeDnahZ3xwimdKVuyEAkvou+rnoWsyhUusi/6Ck10dWENHTSncNMoDet1kdpY3jChJz96M9i4
1ssxP/Z3NB36uTWch0pOzw4v0F8LjhIs2egO3ob1aAGVPJXzjrooQ8dXhNIJu2Y3kKgnBfHATE3N
poezz6+quFAiQD/HVfSba6w/w6gJzVyPlt/D3zhyJJQBU0sif7e8CTfy9G6Bp9JXYwu7D/VynRIN
8+9G4TORVRDCcN9j5ozKhJT8wMrd0iiuP/D2qzPBTMDKKdakWm9Eid4aTMKS632UrQ4LP8Rb/ZSp
JYYRoe6Rv+JDgZp/Reyns688nkRbrRIynvasXj28Ejq84MctGTVNOiOfe/xeaPjRoMghDbZLTKKq
31EhwfhOKNSjVTjDiFP1qBdsXQ2S/gl0S3gwbQLYr0OAr8EuxO/Up7mKVYdOVWtNNGJgIwTWllIL
bCwuP4zpJmKP1Z+9vI+6u+bmIyKBVp4dUVYm6vzjWK9CMP0O7AIivGZc287BGL4NFvjrAyujctcE
4zLWd5P4snjJBnHw7HvOKU6eDucvicYbVnfpW9KPPmqsDWTESCkzicWJZmLpzPYheG15dIMkglF/
vriJcQDvOIDbsdtxUVBw3r4Verb5mCcbLV9u69x8w2xFXQEzhb3qKDc2FzRgc2iBjEgIjJA2SCNC
r/J9NB4jetYrG87dvDyiK9vZac/4mmCx/4k857P+FGtvnIdc7BYmqK/cwMSJ/X7usaueK7XaxrrU
FTKyfCVOH+paX/8Uhwr+Subt4sBVbbhOtCdvu34vKdyb+Mhj2KCV59oBeP3TkHw1WPFoyxTdLcM8
HE7fK9cpLs8YIMEUgTzvZEBfqZNGUMy0+bNdoe3dMeneXcWVGRbHdyqMM9nD8KKmpwzU7VivnLCG
BmwPwIiPS1Sk3aA5S+UR/R6qN/+Z5hNgh2T9J2++n3dAUW7ECGupg7uvJD3OE5UobuyeHR3Tb69R
ANUhMjyJZ0J3fyEQQVUE1npqqVUq3T5lKoTWpfagXIQ12Fy7AdlboXZGvtgIjtwgbOKuq08mOUPd
qDoAbp8OpnHvhfF7YgMfKR5BogGY5t4PRdIMd/ZFf1KtC0+/8MgyKGDjOBp+e7dhsSZja4SsTg6h
82nQ+az74wRh/XKu059lQjGKp0X5FACQxjPHxFxoWMUAa6RigQt8bT3/GPp7HwYWNx8sBFitjnND
9j8isbD5aMnXLraIIVu/RYDT+YdYpKrlYS2sdZtCalzewQrKGT7/830tmrZA/oiqETRsnG/BOviY
ij4MoGfP9POjQ6kwr1wA6y5LKWGCTpuNlFDZBPmd6oGotHDGzQS+ZknyxpPx8vYIJ4g4AT2Xvvb+
Bh4nYQlB7cnWAg82OxT8jQw5LA84C5MYyrcBb2eH5Epz1eGO0b/doaFzVNKn1/tyuVk9GC2OnSAM
/pnggQ7zx5QWgPa9h/wmPitb2mPMBjglgAlsT/TrYhSx1ExnntjWQje+WOtUGFGUEJ34FkgZb0t4
LmIU8+Z2paUmXRDn6QCxzkfK1/hi2vK8yoDqp+Hfh38rKb5lUmejP0Us2Ef+TI021+k6VFDs3eG9
HrPBEjI+kcVH64cRWDvInPxAHx/2lVbC8ELd4uiEOHEHwBYcKw9p2HVBw2fb5L0r9pZbcE9wbEm9
hMUZRkyt55HCTfm8YthzaeE3+VsB17vxa3f7nfYeVDUbdPtrL/sY2hyf8rbiskYITuzq3a2TH4fl
7oOr/qrQJfCjo8u7vqIj0Qs+iNkH/IehauVbH4XfkPFnSEQXNO/+K9AkwbmkLLXtiKSBDeU4NA4A
wjiMfNzrPg4EFl1DfIXPPVlTUEwlZ0z+96CObN9fN0rRsv4FpQ7zfTX2gokB4PZ+Dy4GoNZD6p4l
1RryadHalEvliMehSMeiQvyzBfBsoXNlxKL1DgNl1VRDmN+i+MkKEpS9FS2Lqutjco3JBTDjCmUF
g2hPI2QFtZT/99XVMZ6o0JB1xkBiCobS6pPvZsAFeAwLtPwc2rZjXucooTj5q8d2re5pDuOpXi5f
dx+DtxwfeSCs4F72oS5zIL1smr89bmedfNsa9EOo1p0BhpCHGh35OihMOJA+FU2bjMH4bukhsc8B
PeZ9hHb4lWaWbVgzkMCFOrW/nGe+20GoBBovXuB46mcbhBm3r/Wv1UCqf2wY4EBIzVhtX46UsW20
hEpodZki5U9pD/GaTsK3oeXyDTctd2SR7UIkYSldFeDMGQge/68Lo2zv9CFUJsdyfOu0MY9noV5q
Cl3+5UYo4rnCTCpvYjVw2lnZydr7iVHmbK4PlXi/Q0wlxK9OyVrx2rZOfjITmGVZsidm7UTlPCeF
0aoXl+sw63KIhBwxjEvTGKwxRQV4WeLpkBLfRtDLraEbewE9y0j7cUgkaj9UZ8U3bO09mJHvkahF
l9uJI7DnwRh2PBhsARN2zwJQbAhefjbBr7filmOTeIhXYB3j9rr/FdBeO3UpAhE6ORpKeXhTvptq
QsuNn8kqkrz3FAq5VYIJSi80NlEHWLa8JJgWuJfh/YbjkLfSNlGslUx8LsDoprQgYlEI86nzGpGy
qEijg/k8FnsftD4cna0tQpLudGje7KNJNsnCdWkey1EDkyrrgwOmOBajY6grS3GRZLuCUNoCLbCQ
11CsWA2mng+Khlth9IUAznnv5WVhaVn7PgPETOW9fhPXO5abLAyBOMDD4vOEuem33BP9i1u4eXmB
3AY9vTwrLs1oE9ZoF/eje1uqRxITiRSIjkdD+1FQ47XpFEyZToDAJvjwIkiT2aqB9V6RC4gx5wPj
en1oUtWzQlDfhDJKReWia5kPocljE4JJuYJ0qQMn7eyRrWDLrwAtBX2ew5TQ0TxzavGcDf4E9HQA
Zm5R9evhRuu3h2vTq2agXkJ5zql3Iz+pRecdJDf5YHojlXnrBGqdXGrFeh/GEXl+NgjNIOiTgWt+
hFtX15rMkgT5VDg+YI8OC5KnD7enFXgO/avIQ2gtSa/U5hRsqKf46CW/rfloV/0cVHT96y9nIpQU
s4rHkcXySFTEL01k7cA0Q6UgBXHiH4QTaNzm1++Acd3dTvx/64YlebH64O2GywN0qZ6i9Rk/x/Fd
gCKS6KoZlgULUyfUzUjWcI0U1K7nrEQzWJgVhkP3rDnqsNSxTFrZJTvLmhU+gPBaUft1JFFaIeUo
xX9egaUXTyvLinEKSPTPMN0KZqTV2NwxFechvEfYwyH8eLUslDF7NIBYA5Yn2Gmk618MSHiLKGvK
VflWfCoKBi+GdTUtwXONiqs+i2qOFnbBvTMYO0vArpUl2rfkWr3oAkdznX7prxlqHTuhmjTHIRxc
pe996Xbfpodb4D/RqsA9d9Bb4RAtytn/gVBwTTCKqFsRfzxltQygd9J4rPELopKiXDUsvcpMFVOg
KljMLR9jCCQxsBRmeCanG+P8nb+ZYsTgW7MWivJqs5yG0oOCegKgVD8ppZHs/oM9qDoo170EBucY
KB3Y0t4OLSLIPdVd3mvj/tVQiVgufCt9swFuDZrbHPqZzPJLL/u8Ar3ttkrKh5zvXgeMPEAl6MIj
SoXaul2h+Z3QAUZiCauDgFjDDMyJ9W8yw7zyMIqtgydbUwvT4rtFkK5K/WmrsetXBJ5164lX7ShP
vWEzKRT8dzVpzTTQzZK8UDrxeVxWe2y2Jrj5/+jzcTtn9dlPRBfmQVvfrBvFOFt9bMEJi9sx1ZkM
g2ZW4lFFe9uBdLjiruqLCn+/BfszJzD9czFe4tL69aEn0WUdGqcIQSxioKJEPwuP5SeguucUhX4d
WUpKi5TAQ+GQJYtqZvUaL/vfQBhFYJ1vQ/iWKWMnyec4/BNVke0WH0n20+CSmlnMs5KXxCzuQ6W2
4U1bSXxJt4POkbbYYPmW4UB6+O2hUQOEsYMvRQdOBqpu5H6jLna09cOxme6A8XuKr3E8bj2vtBeT
JuUxhyqefShQ2EJOAr8pP1hxFlx2XBTNdtWKzHZIsY+UQJYrg8GUXqHd66STFErLqIuDvXuUBAa6
EHDSW1v+8HUxf89MWKcmWeAg1smwsZLw6cVUjs9aX/sBX+KXScR2vk5Okb7zOChCG1aJpxesZnw7
BH8LLU2YU0UCj4MAdz9Lt6GEYW4nkJ3XIpew5DzMdiDMLtgeu6pQaQbyI00engMn9vJsNDvEqPeQ
1q8VpsZqhNft1gK/tGNcu01f9wUPG/Vi28BrHQ5M45hH2dy8B+vbtCedjfMm47j9kuKq1p4Zxc5m
PyLOJg2tlVFKxXZqah2QsAZVkgLbmH9LL4vUmxfiyeGn+5Lt3Dhl2H/sRYRuDuRkLqSjDAq59Ou0
3yLsliZtY+gWN4NjOtOFdKrNiq2gtl6ktMl6sfIpy0K/5bVRs1Org0+vFD3mVsTe1tugYRo8vjxC
UUtEsQ9WRQDIlrCkp2ioMpIKo+48GFgmEJfkE2x7KjNfHhDz1LUCCNjdHe5cGTnFqQdTwt0kFJxx
Z/h2r3NpKsq7S3NoYRfOq3fDva9pTsKX7PrDFBgcH6a1oTaW3p83YIVMF9iC7q6sA/3zQt0JJoIA
8EX+BX3vdhFGUyjv481ueIfJm2ail+0ApA17BOMi+/k1kX86ekEXODp6sXK/u3V5UhxR7LsGCL02
BVxBjhTWTLizTjUHySZKn2I8iSenuu2RjOv5s5gR9WaE/hZHFVK/+m9mkYf6do6fRGzR2wF78TEH
v4Niov4WAhXGhqsBRI2a7GrEitU+J4fhIoN2/GU0K5zFbq9qGOAzP4khFJVapT2bfhKWfeVO0MgP
HbN2gyRRIaNaNMkqmODZVJz2BP9G7+Lfd7DfU/6TXc/3/iSkuDkyr8+RM1mn0a+pPuxZh4Wm1lqb
xvV11SNPcKNxjadev3fHS5DFNNgU+e40t1JbzkUtMYh6X61pUWpKu1hYH1AyQ6A+TDW1M0p+YJHG
I2AyW33cvo2uaNnwTwKkl9cp6tzo9PdCeg6NI4vAGt6EFfCS04Q7FZL9wDbABxUKGPlxLB//6QJw
5CVVYcJm3MqOR/dS5PaYVcz1Av3Ww7kNbWb/C8GPqWZofcBDx4ocSWIvyBHatHD0yXkFw6/j2qvh
1p6vmLAPFxvvVvWJI0X+a/eTRWPMt4X3u83ZS8j7n2C9js0hut8e/XAu9D70pcg/ecjhyHdj9A3E
1FMGsvU7yl6QryR56sxRCPuGuESbqLX7GL7vvm5XqEwS7qPLrgQdVUao+c5lDeweYAvs4Zh7AVxP
W50rY14+Edz3Uz2rZfyF1LAvB+cDxs3B0kSw0hKwn1rn7u3Me38hYXw/JsmBKaDYscEVeR8a9VER
Qgu0HRXQEy3YDRYG2bEIoVws/Oq+TvrBzJzgI/30Mw1fJklTZCzznQsw2TFyM+DUJsjyQ15epRDx
B6bqA0EXCufnf++HZZncWDwPPmdFqLysXQKnD4mPaiYaMi0tQELaL49sDNg1BAiSEUP/DYehfHcg
N08YlaDu0O3NtjAQC5D8Irfp/mk76JQjQqRZ5grfME2pMa6PjDekhtPyDjwX2CWpImPp8zunslB5
EAhPE5ORy85mf8tYeLm7bND+AvIuzzM7lskGCuX/t26wi8bd+wiVBBZA+BYEhOiKVdpkiyCfN7Z6
AoWDMTTGm20yn4WpTFYa12v3wdvjcbOILQAXZ5AegCtqrsPzBCHv7lbm7GjsZBW+yheuXUWHsKFs
4wRMQ+jdynsB/OLWrsM734ENXe50Q3vgQfjFQbcqjRijXJXWb4uifykCLkDkMiBfqu52ncHH774Q
XkZlxT4/BkCkBMHQ5zjDn7ZkLDIGij9loC0YsM2hYKHihyYMXYyaqYYygB2hZs8bml8lpK7MUj73
Nxsu2LUS7vLT7P7V/XIqLA5VNzvq4ylqAfbQ3hqGFWuwWM8FQJFTCYf0Lteig4LePfPwRIJcKsCV
/PWpDPdxzXZzTKRWVWXhuqr96TsvhJdCAl/n9AmudnKYUqkG67Jgl0a0mr5Wyze0eli6W9/qeWNB
qsu8S7Pp4nhBVtojmrvohn7QMd6IhNE0JKoCaZoJUalDneG4RtQN4TmH8MPmilAFcate2iBdkJwz
ZspfIv4nDDl9ZB/k4sT+P06OLfJLnwiazRxCav/3qzWMDP+U2/TlAQLbuoU0OQPxB2bc7BV3mYh8
avRFT6eeeU+dvSmKPt/6pORaE9/9hROQnfamf35KyTxNnXKHLT3I5hW0Zm0isKKXJinHZBXLGeWo
XIC/X1/7dqLYwBJxvQXv8E6c3PC9ke6s0MIYZmyX2yxexbGFHg7tHZNZRCEr00qBg3PGDPjMPBmz
jKW7a7/hER5D3VolHodV33l6RNqveUfZG3Q2qMfKUfwNmWtUM27Tbt9X+OZ8YARn1TUje6OGzpQS
ovKPwRUkDMQ1xvB47JRMvRzpN12+EHv9g7bYnSP7Sbq31hXAKCv/Os5fqN0uSfi/zYPeQZMyZDLC
BC6IKg6EVNggj6pXXdLcjIPcA+X6bU8GQBeY78H8QxzSV4PvsKl6ruB+7+sSQCjHzjjGAFZBi9Za
ufY9uWhsDaVFgR07EUOcZ8OeQUD0kgrOU4rfin10iK97A585KpTDXhvGZCCm+/7XVP4+qhM2rVOK
CxqTSM8UGEWfIGwyTktOiRDJoo2TcBIZueRGIKwMYm8GOOhS5+vMZ4ZacPts9KUMPZJOVGJ00+B9
DTr0RDoTH14n31y/9KU/xuF197NoLWG9sh10DYhLZ4AaX63zPK0eKSPWSTunrku2mRRKH4+np/WK
CcA/kTJsm2KzIOhSTCYMOxSS08q+jwkpnI35DthjiEdQTFjnCsRQsQH06TyAA8K8tNwazo1kEoOl
Qz2t3lzv8EM3yCrDysxQLk3gMENXzsuUKYd7VfbrwaxHefmjoqm4Vzzo4ciwIIky+VKiBLrfJeln
M9xwF+DJRnhRS+LCe/oxXnKWNCzDWP+yApKbQLcusJuDHxGy8b6993S9FlNZRY3JRlqtt0A97c68
bty71y/dSxGf/ciA6BSkq4KjuRkg954r/kkco4sUXB/LE4DETOOZ1ntMK9q4d+lKlabZEucDsJNV
MOh+usXPf40uhJTKt14GJW9KHEHVWzigLGt9pzrA3Z9jUt4nAmheufbHRKtXnD0kipLNK9ZUgbbZ
nCBtEpr15JRYM24Pis5qLJEGYzCPm6Rs04+JoWlesU7vwltK00EuVnpHSxDfrolMWSjmrLID4s5I
fJDbZEjgQC3NvKThDZxitlCJWaf9yniDRZyyajd8qetYgzzCoHt2nn7tl22/ivV3OM/MrFUTazpi
rQIzHORaW6k7r1QsOdnbkyRq5gqG5PupUg4rSLkVLAMWzbRF4anbVhkpnnj/to+6FrMY8smRTG4M
TnHFG/rmassbYNCGaGR9fHvu8S0+zh+WhraonsvjmJqym6QDF8YGdo9S1VOdEGh/DlCg6PrikkkX
dBpcQLW7L2+NRECavxUz0uzYG65Y0XlK2tMNLMqslYNIFcF4ZNHHPizoD0EXX7LSL1M2Dv86MiMp
Uo1ASZ696yuVAUYFDrXWOcQpGKRHG8I9BnhX34AC3LTJlL/HUuxe2kzW6ZXmGtxA8OHs6RAHgKQs
jqqTFThRXSz+xYYV4RURudCrAUT/kKwGTeVEHg/9lCUBi1xevQ+wgj/S3hHcLsgRBl72HP1D32Gw
29AMxkfPTgx6hlQ/CPz3+1MtX02ENY3AlFhQJDgtuDnhXOzFmozO1rCa/fRcmrdOBjlFnk+tTG1w
Df9DBl213Q0YIS091nDPXAFyB5D7anb6MMHDs9htMQH4aJ1i/V9kJFd61P5hadDKJcY7ubkCYIWF
a2pmJEOFYDRVbyUKhD0q3c0KSoeDxzqCCg/WVkb5bA3G/NqCbQIwtIVeTyqxfK00FNIZ7z3pR1vW
+ZCbaBnA/pV+tvZw296r0inWhtsPHUTX0DoaQeoXUgPFa7m+fCuY/awanS/WAX855Gsyu0ZVDWso
Kf3u5TrAYAXOa0TQCyvhwZpV1m9d+HWNxtEewg4Fe7pz2dfyyfmmXiiLX17NQNH5Sb9hGBibRrrK
/vwdTP39d9Uk5biNDvaKEvo+90iGEf9gmFnY757ixvKCBMCDxzWQVvmrouci1+09sGsgbm62TucG
T/qlHCsuDzKln/NcI9ksl2sY4ezKCjb/SE4U+CEq8Q5WbHJFiLuvigo/3N0l/MRWoNlkYax2QzVV
KE10XUCkv5SrJn+6inF255T9mDhS5NIYaMRn18qoTt2jl2my4JAth/2lYU3xt40924Tbg7WLKiOZ
1pRXOY3j2ZwtvJn0VRCUCQIKbX7yQqVBArE0EaaX8vBgXMXMxQYXL9Sf7gKOrXBY9kjNZIAR1RGu
Tc46VfUAqhQIof58FA2tgRM13LX8p1cCq6BPmMffHS57ARV56i7+RP8W1NxeF7snQfVUN7LB99tT
nTBchn1y9h74ODN47cxcx6TalTxkijFl8F0yscuLnUd8OirjBl/btQAzKY/Gg2TZHHuWjqewoxk6
52cLR84PDksjsoxooAHba1GMkwRT/AtQ1CYS7IdpxKBm0+bpR66hyCUEmLNPLVeF4IIBA+B2gTRa
YxC9jp3wFE9pU6Wv8THKZa2frDe/NcHir2J01sa5BXaytqoGXicmdhatHDNtw7bVpOQea98Ma4gF
qet8e1AhrxTRLnMLPGDWdZuPe/KySmiyfId199X8jkyPRz2hHTce3MOb29sDrzqlWUvAPQbBBFQB
X+1Bg9NqB57lMidaw/ThAlSVTi0Sy6tgyrLxPU2bxd15MFNkDcPGwTlkmga2Ok2nniOcG2/TsUUp
fkVQJcFPiX0UWBoUTBWG7Djl/swOGI3f7CP0HnADahiEYGC2JGNYnLcOHMBzAEzJGV2ajvlW5dA6
El7s1sFVV1QWmakeYnVt6Qrk8S5RqGvExwa2a316wSCYGn1SX2fCyc1pHlwFRWiVI29J8xt//qfR
54m/RCBscSR2pjBMHTl8z+3AVYldu9SOpXs0Lok/yM5gFDIQ5RLZw29n+D2vyJBFy/ai09YleEoS
kKOJqwyaSEeYj8Y+I8l+hhOtF8B6i4LcaBbVhGYplYnCSnwjpLhGWy0SJkYP9JM17C3jfqubpss2
MqH/VW+SUY+LmP53TrpM2AhYPJW5ML4pvXv1/Mb3+XgaZYu7rxnB3di52D128oSd+xK9R0jWWZBt
93mOTJQm8FnzdOCS+8tl86c2A2RIFBrhPxE/wllzj2AOI+L71usScxLgHEZPXhfE8jg8EiKVgEeb
Ez853lD/QlcupIIhb6RQZQvHOodOBTmy9YN8NPjbCb6RPJ0ZKG+1G2y5GepfhbZq9G/qLyxLKe5m
/ii29+NuZUwPtteWqVFN4+46I1O9ncDShHTMeKXejEt3kKi/n2Q9qR/zv/9z3xhpiIAGDdHaf9Fi
V1u2Blrf/cHwmM7IkwCju1kXNnfvHNZC4IsqwN3b5YEggDzJIB2Qqs5Hr7TBpI/Amm86bT1vfb0F
L/pfdfZw43/OS4XTDXoWwamPgIQa4kV/+CCz/VnAB3GxDCFH6l71SaRMStsHSO9DwzETYHzceivN
pSfqW0EWft2uqSqTtLHEVTURXSma0iEkJyHoB6C5j1tZ1yegoMFqMCO4V8sissw8ZvtLpc23FTSs
W5O121xantFtLqJ0ISmgta0pBH9onm0Oz6sfUJGu0pIEjHA3+oiJUTQmlgJscLm5eEbkFR+M7++7
Xq5lqB/c2P+tM1HcP1aPcjfp1XOO0eoabb9pc6uM5LeLTtPWHRPkdPjVgNFMdi3Er2m3SoazWYYi
34fF6rUoT891FrXSv7weP8jXMDG/EqAmt87gSmEJFcGRXeOO80RsSJlJCV02YcvA4UkL4RIZVR4l
KCbPvpfakaP0sembGjC8meB5IJhGjR/fdbYVfCTBk0Lr9Ijj0TGDoEtfntgALKy5RuEgb9pVWFoT
N7+b0BRIeqPcOg3mvP3ERkYmPf3u2VYpvEjUvvvxPEPf5KcvLLnFeo/uegD35MbQX2xYnuHQcsvz
asreGB1Ufla4w9hVNZqs5gwJ5Fvl2FmQtiaqLXRoR7BRfxURzXT3NAeJouXNILcvWA+/L3jkT7+t
cJ06pdiYytIlyZQuPVx9MlwV1ctQ98ow7nhDWB+kT/xCCQELfzZo2q1s/tvGxxooIiOzMUYQwD4y
mGmKY8zunMPqhpnOKJyNWCkgv7GaRsG2aH3/Ss1HwfJ/pa4Q1BOcUjd1aSrdYZD0tQBOSvaAWvgG
INAgfIPdZpYkSy33xk6/fNqHCRU45HpdbNKuxNJ3Ul2t79tYgWEX0pa5xoQjip+V/+aBk4ZRieoX
gwqIc5U2nKo5v6u/uFL5f3KTX2pR/Xvl7OhaoglN/f9FF1b8sYdBq0kOxIhruf56JBTRtldr6MeN
NDS5RwrbbbuLRTqGxtwrHViAnRbKkfp635k5k0hq3KMDozkiDSmRjLjYgM2ZqZT3C8rGoDR6q9e1
vZk6+NLEyxLuiybQcYyvDtn+vH665OAQqBm91XMgw0+uebWBmRYtzjO8EVo9JUYWTDLGgcaHl974
CsU2EEu+YtbyF9JFMKxCN9N2rz8hTpPsXNYAjdQO65N5NQUKyB/RjBTP3NVurm2XGigsOdf6O+y5
zFtg4Fn1eM/6a5ul7GiT1vtLBusPRKuV/kGqxUIU2myKx3Bh0uEEKiuC4a4D3YLHhEL9rKmMQm/P
5qiWGyvk/svbanBXhTikqUD9d7kXs7ziWPQaWpDQ7CikPCL5P666CncTZYwtfMl6xn9NygKZ7Tgx
FQ7T4z0YaVxlqPtSarDySuasooIABebuI+uQh7WEGjEySghq1tMXe6puvUIVe/3AEpPWk5ZnJF+w
Dc4kQpBMv6mmhhjHVGeDuZ4Q8ViU4rH1cxkcCpoms5Yp2Uo7/B2WxeJtLaQ/GwYghKjovwrRua3k
k8EwlH4sJGgKaoByip8Os5c9ubfCGvU2LJoTEAhLu8JLfhcfdI098mt24BReECpI1fWK4Tzjvx4L
aUaduLdiydkkKhtO07dO+7NUAt0FwC47mSsXgZ/VJ7BDR/mVQIetHmBYF+V/m+HAf9EclARF6TY4
AWOx+uqrbw/kUIGmDzK6xK2hcscZLNnV9hXUMwMGKk2CTiX6kjj6hzWZ4dvLXywzmb1xic0DWeQt
wza5jz47+dRV+WlxYlYoWVtw+Jk9w0b12i2lSEkYUoyZpk/kWi7Sa0/hL2ajjrXtUhql8LsUbwaW
BmGEEbH5AsPyA1cQETDPpUZ8ACnIvQtr+WDD56ky+I7jr6qWAfvK/vBpvSkCB3U7SAn/+L/H0WtF
ZRXkPA1GdjDtmoB7dF8DQLib/271fWXkaIo7AfnEp6t9iCgyJOOTpi99VZETW6UbLAx32cycPPXO
t4sL/DqvzuDkAsF8UAFEfHUT/v8dl2i8s7rC
`protect end_protected
