`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EvXlztZuzLdu/k/gvCmwT3YNPgnirLbxu8t9LRgszVr1smXiC+eGAtTIy2xF1RwPiBjQ7ywg2zDn
RBc3OAdot4SiMpnZHdvp4iSUeU8IRGBCV6fFvzkljz62wLVnEeVvVKBV6EK9weqxPBbsSXriosA7
JIT9P/8qFVvTsv0kfRAf6HRtJj5o2evFrK5SzqKnT11yNQGz8r869CbXHF+HPL7DUlVKgH9JEV8V
7AW3an2f0+cs3cGuSvjJMZNgRvMnHgu6ZUXlH9bjvh2yvhvFzMZ6Kjjem1/+AWdESKVkoYi43K5q
ZnQjZZLnd1CYh+cHoPC/pG053mgikaGgL+k55g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16224)
`protect data_block
tMmXiq8JZZM3EIUyu0UBzI79amew1gM126gdrG1H6IJiv4UfW9u41fR1BczAs5Vv7u2vUp/ND9K4
5b0oRH86KSVxHBGmTUhYoNN03hibHpR5b2HD31NSQO7c35BgjJibMz+Bkeus7Kp2Jb2FG+y/HROj
XTqpRDM0wIkvl2cAWibSbBKyPnVDk5chZFcwxmMPTmgLvId7m3vsgmVZFcBT3EKxX0YOeHdb6nAu
S1MX+yzbK+0qUrtOfCo+HtjKavrIsM4/jKrKCP+CdrSqn3+JJqeDZDYvvW/YR09+X43yjOQAsCnw
NBsozYHMjDKliZsF713VG8YKtGywBPJcx+Ttp8XqcOKK6AIVkbJIaxIXJnDfV0benp1eyPjQmSYs
HJjyF3MhYwubZeCGENDzPwTzTaFLB98AxjTIudy4l2fpoea/CbY6LpR4SMQJ0GLw9lg/wdb5fayJ
4wHqc+jidz3GvOhG/ycjgJFjtkV7NFQS79JcK6KCtSxoSNVWNSnbF1uck/mE1mfK+4H+qS3AFSoA
XKUQt0aAi2t5up4Beh0ERx0A8tNeFKgXg0dL2W5JJWva65ptpF/4vBApBbq9Xh3xheM4lPCi4zOd
Wjgmc/5JGHKyQ4dCXKp9ktZqI6IK3dhqv/gvQLyIxa14uSUa0sxrimlwfAmBP5k542uy1BXNXN+t
6GrEPESZxVLzcj+sdMGF2igmWQwVVJ3M2+wl8emTFNTYXyvQ7DG9S4cz4/WgJiuG9vzFsf/alv+W
LWrRlK8Gb6t1GMbq2u7ZXKGF1dES0ru2LGC5W+nfSF6/kx3be1eRWli2gAAa97xvTC+LO4+KRrVt
zb1yNwt+PUZtV+KTE3/kG7yrsNhiEPEPvmXfHDG3i7xDUSmIvdHFAyWSMVUc8wxxoXEejlD0jPF5
BL0AAX6ufzhfeJE3mrUzE87HhHnlbtux7k4a/OV4K5EsySuGlGrODqUWxURFizolj/1n7kEtQin7
BHgx26/tV1mr2kPVPQY1b2UqIjuo0QwTnl/ZILeOPnI33MSMMYaoXQQyxyf33yPRWoPdjAWPb8mW
wDGovMYJ5DRU8fS4seDrNWJHMUWe/VesBOKNEEvhCfb05RwoUWXUjwW6Ij/s3nBFvPcJOeule0vI
Q+TVYLxo+GdIpy3Jw0CnnpzqEc7dz5tGRL/Q2G76v3eqVlzCavFJOYGLA5de//Z6/DjAgJ26kP/0
6cx9oC497n9z+3VhWN5DjWKp/4xpkgbK3QMNizMygrJibEiOM0BhJM55ZO8SteEsXSf5C6744w89
GHfuAVL7p6FJz73/A7XboaF5gYD/F3FpKDSBTA/NrnD4hVpDdAijRAYDJHqfkBG1OC5+HTFlzPQ4
Jdi7BD7LaebRjYEG9DQ+UtTWecophnbdKDQVWDhezGfW/KQzpQKL5zdtIrbebeQq2IATNaLRJVbT
RAFoL/491AHwZGHt09NhyxF8qV1d/tZV+Byn0nvdCJd+6eStHl8VSejlw+1I7jOJFvH7ONtxVfTM
kCwQVko+x968oYEES8X+xXCAUOsapUULoukY0EmJeNeFyULVNc4GTuxtQ5Hjhc6ocLMddles+2Vg
tHvkDo2g4qLyaniqP60FnvsG7eJYBJW/CRHHHSWNkJSc7B/RwTDZNv4XHAO6XTCMeBsHFIYPdz6j
TUk2k6/ClGkJxhCMM0pDRmTJIVn8yLQhws3W28YjFTYqGE22dWApACQrziIoXWytxnBunrgwQl3S
GxK8yUjYZCGbFimEmKXe2Y4wMm/+LQ/IXfJAUE6YiXTQElj5Si3yjkecuHJ530bFFlRHzfLtuCc1
xDPoDdMNfXsZnDUokqh7yYi4uqepkEM1EIjkek5xG+WF4O+Z0LdqvtBpqGLHotoT5kAPm47rzy8/
KA5voR/0EyuUpWpbB0ZR7fHV9uzXbg8ybGlwzxxecdajEcWeI5dQVyZNA0sqwolF4zL9ARSCsB2t
cjPya/45yeGb4vFNsZ4OMJFtgXi3JCvCg3g4z00MgO80QJFyrzGVhEheHln6cb12sQ8nN6yq9kfi
4+nACygS+O9EEwow4ZK2jUkyFvjdJniY1psyaKq77HhNMwrTQ6vjzEmGIP/QScqzej4jpCCDKfbz
8RhVZfVM9rRG3XS1Hwz7OnRB1XPLU7MDw49wKK6efI39hS9pegpO7rletaKxI4BRmVkCBqOgPzTq
Njs+1LstLEJ7Ahici5T+ZbAV8+c9dtEzNPdSbku2iug3Sh5S86un47TAdhGUboS/wCy3mrEXCcvN
wPfvzb0E3ed8j6ZdSHB+DSWj0zrs9TptoueyKrkBs/tixIOkSNbCZvO8sv3TI8ZnN5BLahAXI/b7
OUpEvE2ZDD8uqu7ee+J5OXv2sY0SsRV8b3Q1mDwkfhVRwU4GCsk0H/foy6XcwOTp2NmbXhVcYjO6
+bllh+iq5Q0rT7/a/Za0YDRXAYZGlkJSh48YFBE6WjXCMylSvcQflLLR3aVinma5MHG4OUVYgHMO
le/3iY/jT0AaTRdCR/S13fq+W5r0/dTYCit1lbJG7FCWE7rbHd79+aScTxFdLtMINaL4x/AxL7R5
krsqcaB0qCvplxcyLjCqmSvv5XsdEBaVuMUm6r9lXGxVC6M7skxfAFUmj/FhV2H0PWnBHbfbRD0w
GIWjpuO77mSOSJSFab7TurgKAwmWgWIQ3xMxAf1Gpzf9Udlmtb8InJ+6ZEpi2RH3c6wr6zs5/8GZ
qvaHsbpijTRTls6XIrwD7UPbiXL6WysNHX/fRZgfCMT6fKf764xXr9T1BQUxcHmk3ywuX+z3u00T
F1TTmaPFnaNO9q0LUqrdE4e4qNxJqWLzzQizjRWK99Kns+6pVwcLuHpfxexsBsEAglrfsZB/BBLW
rOREwRY0GANQZplu6zRDDoG7MLReFQzlkTtmY3VTHkpSyAy5E4KUykG9xLdMSDdO5vRHss7Z2IOX
LDPkqbVxg7cnMHrGsrjzdXTbkysTSm6s7rXaKdZpjAK8mYg6X8joAjpuXX/oDmQrbMI35acC2lqS
aL8Gy+05vTT00P4i1n3gw9K/WX5CzDtyyPniPt2HEA2i8OWnS/WyfUHJq5vQ21xb/dFYLC/trVq7
fGWV3xJDlcuXrNyIXwMXL5e00b1zZhURE9wJdSY6SSb//Va3zBOSTv19PnfcE06aX9taLCJ53fsd
hWWcunyCj/qvE0s8bIgDOwVjcMJO3rzeTP3ETT+xG8/AdDx2HdiCY5IwAO5LoPD7nOyqqz6CIB/w
+AnyCEQeI9xZJA8UmMof0WZ2AMpVXB0WRE2cLe6KCjlmeKzHw6FYXR+TgwPJwAJgbbCbEqEYqRST
FmBJXJSBsqp3t6bOFZq84zkV5zuMDLU+XW8H9ygSNwlmEe7CJHjdQv8I3ahAz1J7KFwzD+UB3q+2
wm9/2F6+++YSvvq7y5T0McvfJrRN/IEhZHLg9UUxgHFawEEqdqCydUG3lSecgObwimyDFOvzKcby
QYeVlG+RwgRNRpWWZoy3MbLSNpXZIJ9JUz9zd4mx5Bj7063wOY2x4XOxCTo7dfUsxi55hi/GQyZy
ttC+LPjp6483A/Z61cCc/Tio3mw6nvymAtZ3scn1SPdZpTOrQeUGbCKgSq+bZluc4zwBg20Syx5i
84lnjrtg4rSft22g0d9TVBNrZ9+KiAWfruqeSmBkroRvwNiTGoDRGpwEw0uvejK2NkM7jZkAKaDM
F4/pUpiHbWQE8JWbAtRb95A+IDWvCgsmPV4msT64f/N86vMfmwNtShovbzmnmXewHxUydGZciFVh
w6tUnlMmiEnHtRZLTMQbOwaF9fN0COGIlhE9GWMiBbJoGE6i+FSNLZECDa3ZckDT/L0h+DkFFNmc
C43jO8YkS7o+TpzmM9nNaUvySZ4wnuvaX3W6Ibe38qAvML7rS9hZ7/5OS0+JRzqgOs+V6DpstRG/
pwsWMCZ31LVPhRnUpUKql1A24YfjqZhJMrT5Z4rAoLB2kHVvXAO3RGVaEEv3iXipFE9L3kSzF3Yf
8LsoPEHN3mDuZIRHiVF3MsGxg8SkuJ0w6LHDGtcd+bqIlisFIDZtR8r5I/umlHiGGKA2tenRoxvm
gkH8nX5VM9KcKAqb9Bn8I84VoyWLu5zYOSKeTbn2qly/CgoRuHHPb+dIXer/Hjkc+lzgfIm7nneq
cBvO1UMvRczjvpoMg4D11isGakwwt176Qwq9RWBU0S5zuR/fsKlo+CONU22O+XSSsV+fYX+nGI/X
syosZ3YewBGgiQlp+xmb3i+7Tj4xa5BxeXyWqfh4f2FuEgdTf19UfzgQnGd/d+rQvFz7UN851C6m
Jz6AHM2JsgOCuvV+d2TwAz2a/GE+dncOMv+HgcCR6ToLDJnSsIeXAzx06H2eFdiKzNJuHHjGvQIm
l0j5YDQ9xIW8y/9fOG54cPPCOHLoMn7V1UOLT7dfWJo8JvFHK3l5lvx+0TGA3Na4PDgL6J3Kphn1
ehSz7M7cP4fb5aW25z80iViC5YX2RsCzYfrfZTj110I0dFlBIu604hPHyy0vg8tDonjMUJ1WI+sC
bdLsj0N5QWcEkZJ56bDgOcnqHp43gUNo2gr1/AwQlkG8lcKlUVx9wSL48CY5fszWtuLGzJ4JVMnL
3D1ryX36MjM5TIMhg9PZ+pekTGoo+2a5tMFw+t0I6NDTzsxgK6eorBFsBQxSGs4mwh5XWxIVLP77
1FMqFkY3vNucEzWthbrsFJ8lfj4TOxZd9Wuc0qHn1HS2FU9NCLj5fjT/AZumXAwpf1ENQdeot4SQ
htFzkSEXhBMRgecYYV1VPzKbcfVdgpa1WSEigV4bC9FYwu7KH8Lck4jGpv4XdBnwRx9cDudlNXpO
9YkbRiKuxkHq68u4uY7Gi4IOej0JSC0TotTpwRfT1BUg72HS7LSreKJnenIePoEsn4HNjRnqBiWg
SVU9g3fybVXYhMi2968XDeZQGQNjE2gKWZ7Ubs+koHDhkEosDdW5JNAr4KUi7Fnm0Q7wSxw6EP8L
rJXieMPSNU8/ffskFtqeVdDyNyu0pGGKjiVmdog7MytFwt6ASwJO/wvmh6qHx6pvxRkCac/WLgXK
wO4q2Wf2bCdqBp02G2/h+C2SoH+k5FVxnN7EIgrVjGE4e3PTstKsD9Pxkkvd+6ts44sfQ2oWEi30
hz46S8XSpiAV7ibhkug+gv2/dwM/lInCWOozYpXmYgc8+9b+sKdAc978FN2C0ZekQvJam43+uiUU
VZzO6qqgdbnfWX7kOx2CbmtdhJP3wS/6h3VxP38ujEh6BkqqtOeZw1BekyOUL5IOHo9H45yv4Bhw
M0nj3I7WVrQrAhlkgDyHVRoWaTp0rXKO0SJ6JoGHOn7atN3BkXG995yPi93uOiZ+XPyOyV6+DRqY
F8B8J968QBnE8Mk4wRTZaE0/B0I5Jx3RHUDfC8H+cOaZQKLszAbtA8PkfMM/2t/m0TwPwO6D9D7d
sqeKsStxicCm6PNp9hg1m60MAeU1Q/7ch0NNx6eSP3UUFBMQVnXGV287le1VaVNz0Dm+lK9s+AiS
MNNRur7uJit7YBeM1IVqN1aZLrUDuNNJJUV40WZgj+BtQ+JKh2DtXunVJ7YPUNu+2QXMPoyhtc25
QVPAuHHe4ujPJgmbBlxCamQkZs/bKhiGzTBO6bsptggdwYRqgHUW/+uaqb+SXh0Idgm84KKTozP7
yBxzsiqNEhBgqe0jg2fkziVwDK0IKxmkubW7G/XSMH7fDbH7mldLMmK29RaHXTv1NmNtxWmEubEL
msvGbzIDw8giMm9HjYfC+mqaCBnOEQ/XdsFZsTeyeMim35eO9JQBK+aHh3zBRcssoxeF1bcoaco+
j60GFLl7Yn/6Z9THBT04XPBxL/ySHy254XRUn77zt+0gR/93rWNYoVH0rQRrgveozVgJ1uBMFPUE
laIMz7jajynbGoFnZeqWg7jPBx4SiBQpO44akaLXdlKuH/XeVwCWe9Z7D0PiJrHyGH3Z4hedovjf
d+VlDduwRq7YhTufy9RAKw2xuMSuYXKQTPmRGjuGo5vagr8BKQScyuLBg2RSEBMK6cRm/05XMXAE
7/gVeCGdGvBZhUd+z9YhtSP8Cj/RPtVIbvM1LEIfHz1DjB1VucX2vkr4Y+wBbyFvqs6cQKD8gNUG
Ph2fHTjJah23cCyCu4pmcjEJ0tao/mj3eEQ3a8iaVo8t76NnLxqQC6+nXZoW5A0J5IkWXqZBRfMm
ZoF1MHEnWef5VzXXwqMpmWY2N1RkFHsdHT5vTFzrIFOv1sjYK8fPl6OobPMKBsNqstmb9AuWf/Wu
TCnYVp82e4OZWWuL/KkmiFRwLuJhgC6HLowa9UhrsjcA2rHVTUDZokpBySjAIFuqi+IfO5/mPZaj
gHiOtEnHy0SlPDRn06yMHM9Ec1MQKKZmi6dxzW4Lk+F4b7fxiP8Sg1hMF4nJHHYAv18NP/yRq7tC
NoAK2jFOrBWuiuNgFS4t/QeYmJyn+bs4QPr4ikJjkP7Zsvf4ipCBUuW8JjOkeSc7BwryP5EZ14TA
lGqC3Pdkn8ztubMq5uS+6WxmuuGfjrGXcPQpxlR8g98FwCcod+MIv3NRwm77cMz4R8wdxaUTUCit
Gp7IGSv3a7W9sWyp8ZM+5GjjcDJuR6AMjXvrGV54H18Sx4kanmaVhwVNW3KmMB57F+4I2/a73LiL
3N0rNlPHQfYtXZ8MdhkTMZZoNG56npnWp0+pFvKKHJWk0oyYXpc6B2SHdL7eZ4WbjYV4FoSPH9ac
b5LXxHde/8Bfl8jyo3u4Q9cDjpJMYIEQH4LkGhpkFb9TsJ+/0z3ggAyhu6amxP9PT5Ps0SX7LOTA
c9KpbPJtRxquUqOh9utUEQlpMlljevlxBHX6SWyr1UpQWfz/rT4NUjCZEf/UQG9qZV2VMdqVlhep
U0Yd8OVKbuiLskr7oU6MKoeSqc7EtNhJqGhurAP2Y+4V2+IrO0BFv1W9KJsoakZZ+9aJND76/sdJ
1o75ciVnL/CqHkn8vuzxBD34n4KjeuB0g6u5H28dcMaQqK2mTEdGNoY2dH/Pck5CRmVjaNb7D+gq
8LuodSLjv34Q66cojMmiXUblSUegSyceShdPIgbMJ1Ckonn8uNYhTEV6VKL8fflxzFtHNOYBBXpt
M4HI2Xfe4fysTVuGD4G5/Ft1AygCjxAXi2zs+iuMwUjjiSjLt2dEx/zVVgYR4jsq/wv0ym/JPz1z
0w60eEvHWTuWFhe9417PnO54ec5u5OGEgkqYaU55TUarVwY2epRPbKZIR00OFtawN7Q1Wd7I8fwH
NZPg67y5NCgJJXMdjD/R/T+bSFP1QdL2+l59sPxNd9oxV+DnuJjPTYSho/ujU0/S7d1KZhPvJ0TX
PRB3HIPHyPoCIuf2lEzJ+AqRNBVP/z92zT72QHpkwqQwJHJSPHZgtDsUGK5ZBUFgN9mp8P2LeYPV
fH/2lmVqtNA9taIKOLkX6ZJLW7zZUCGT+QPPUYvt20E8eqQwVGX7/SEi5c+3+hM6u2kr8A6hQ/Hj
uh05v+4g564dkssO0AJCJSEGruJR9XAc0kt60zoDI8ZfPC8/ZCC0ZWNYu4EoeaEBqJ9Ez4jYKBjp
7q7Yh0wqpKfyZo3vjnTgftaCYEry0/cKNIB88ffrjoO3X7Aepyk3iJHBxf9zUdt+x6psBreQyA62
YMLBsEBoTjd+WIg+BgagtFoJcfAc3j5XweQ8zCesurFAbbkBaABuHouj8v7vrKUd7210tADxBf/W
K5N4W2fr4GdtxH+rGmwjXpCn22JLz7bFTvmYAMJsIWe4Xa87UB9KHzzcQJspXuqXwJaZOKN2rkok
ablARw6dgqELNcDLvpc8XjNlOpUwKDwLG6J8FeQv85eFL31f3Rws33RNPo2luJpk/oK9Y6Kx0QY+
U5pKiTR455LfVse1UcGKS7g/UYxEkvEoEuesmLFUSNpddjkbTvYMo4omkXHmM6RuyfK3EwclWYak
MCyld2SFx/n3bIoq01hEszE1iVxaVmf2RgRYCg/aBdrwzTrD4qfvZp4D1u4GCVGquUid4C4LiCRq
5E/f8Snf4G3L1JaCeVg7mzOS6J12/ZYg961BDKTUizJQpaED5e0LdzWPDXF+2RjOzrGsRxPDfd4l
QYtibOnoB70ogICtOtRxLjHQoMdaLZodaxFsxtTDGmwT8GoFBCb5COnImxeCwJZd2+SlQOMzagj1
d0NqhnnFPiagqI2kiRiJvaJDHRVsnNPETBhqKjvrouPZDidSaDA8poNYq98o5BOQpKkKna86aLPo
n7MPgZIP8L8SarQC9gFuQos6dhl4QgpgkBtvzfkVHAinycSb6/Vxs8yY2A0+0qg6kPcXdudaYUnY
Awo9vrCCtfwsgspzDNgb0DQ45x074ZZfFk7zlXLQOoWTuUWiCwlUaEa29Y3s7B5Gdl6oNkA1Y1sr
xiIGOf3tpdGn8EGZJ2OE0W18ilsARDchMAtuvndDzmPb8GZWWyOaa6qJB42FaCVWzV42msHPiR1E
IawA8LdgbjbMPk59llJGa9CFkKlUHcSeIU4AShAJpzLneKxCuidXB7fCdaA9/2G/2iwyLaVkj4mm
nsuzwn5syPWEI4CM6CAQSZM6APiv/EA1m5AvB8Dq2hlfYonEUKe1W6gYkvmXMgGcKEY81AuHe74P
vdjvnnZuhHINuMG3xsh3mQblmbINSHSc+GKKcLqLnquQ/kMwy/fIluJZoTyMGvM0mKnOX/YNlLtp
1PIo457XgpWoOBE5wOz0ppNUQuN6RoMAQDZUnqPwY6CPlEkH0AiyowDJidkzZfLIhRwL5DEBmRdA
T7oEgpsahk9m9QN+JLQnvmy47P8xG7US7Nyx5mmE2MXzQ72Nlq8EygvHacUADwfG6Efm/+IlgPMP
S2m2AZr4dYpQMp9+hWCEySzyFWXm8QX5YUBcrfXzrm2DqgsP8yvrwD92uRz95cmQ+GtbPVZbZh0X
x0uw/2K9gleTIryL4DIZg8S2bkwpDiZjfqdPI5GcoPLjip2ZCNFgnCNZGYwCgawzR64Bai+9DvD+
vBnQvTq3M217c2G26uYoZY4yNk/Ch1LY00yTJOt/4YYJzayvPT+m7LKvB/+UCLpFmsz1ED3b/wRB
rlz0c75LLw5lJCV5xW7gsKZaRdJMaTzAs2vOpbLPvdhELT0IARQTJp/TApwNiWiA5NORIhHQPRoQ
JLYOSzYCFcPmtISfxVSjEV6ecu7b2mXt/RwCUVNlfTrgWQZno74ZY5D35zFlmgcvW1abT/YAfw/k
KMiVC6GWgolKvZ27V8ytpU/g+YKg2hnzZF6SFi/SERvQyuTp59jPzRK6D9d45gn7GDExjujtSL+E
jXC6VlugPexJy+WU2irB2d6n/M4XHB1e6xiaPOpcylzFWxQ7QIL5ZWjIK2K+I1ZzhB3H8Rwdvqqz
ntSWnldspTrdVT4exsn2HhNYyBcl96c3UBjpmLpug2o/wqT9QRDVqvkI3ykEGqNxoCRvom1hwjck
fAKdhlsmXnVdoWE1zkRIG7hEMHw7XiE6JHVhJmz35vCovoDF9NJ9A9d/DIx2uEgAjvvAKABwZPYp
Dph2PmtanzqcK3mkMNQzxvxLkLxeNtVsaQL4Y8GQrlLzmOExnTBPnBEgMMhHi5BRDUv7CdN5NOg4
n6xdPwDfSPoilWr69BUA+iAvLvuYKOs+HD/MzUCb/aPyAm5WOnkUXRzC7F6osptZldp51+LgePVa
BNsv5TD8Ju1Xt/TAyaoEWfERiJnPhJ78BOHIyV8amNCAE0vy3O03+Fr9cRUlAUrndW/WzVZZ90F4
SfXC2zDxo9mYHQkvRAbuohIM6oqiTo3Rav1fgHgywU3F82T0JQ9IYnslGfAdRGRdsoe2ertvV8g9
oLoOXoL5BnJhfG22mGwGmF5BYdxqX6ELxt4+/RSbX9vmie/hVdgZ0LEvD3Ocdet4nGtg4xUyq1A8
PNRmC827dxSvTy9uo23phrWIUwjPEHjuevuEvjX/sHljcAt8LE5qxHTzf34ZfEfLjXrEvLWNC3lE
cPXTNhD4akwHj3bISL8mqjd/J/uGPsJk2+D0sN8JTKOKEI2N3t3TQrKULxcAuhYIvBdmLwsja3qx
ydZXnk1GTbDEpjwhfv12Tk3hUu2ZFggEzG6jg0hH7kyG6LrAM/Md1WzhbMHs7scvds+w+HxhtgWk
QsUnCq/djOQ1m8KLhvvnFpSuYfrGONBRxYT2620CLGJHHQTXLMHzNERrEPXFaBxs4UW5UOxvRlFy
VEuWZAEatp1WI0st1Ez7EAkgippPIhd44/tkpiRZDUlCR4uhA+PQkV60XEpxda9/5qvid7XuG0JF
wmTBBscQ4p8eXU8fc2dJ9/CS3JT+aMLlWIgCnvI9iH2WbVd0W45GfNuCcH3o9YYpaXcmjr9cKj8C
4dovrkyo5cyy+7DTWYSwO3CJpeSDIH2FmWrUin4pZgHMh+C4avz5NuLDvv0rne/CM/ZBCo4QXwTM
lFsB76ZiQRTLW2WNSy6LaP1J6wSYPikQHpkS8gsPj/mn0lXExqkW2x/nfySHAFQXLnFr/ydTAE9k
eTDh65McK7NWq0KCs4yb/Zs6z4Hz0efOeu96ecCm2VAZnUpzUS9LX4Q8SSl/BHyWaYQbIlzr1fS1
6EYqFQhD5OhUer8xa97sUBf1mQK4WKpkCQsAIag5hhLwjxkHNvJI+TNH9io0sWdStHBd4F0L/GV/
hufM+3jr0arndQQXv0o3+9cXDgqsX01LAIvMJYp8XvQeD2d+khh+rufYGyZwt82y/pH1fJ99Iryo
91tDVkYvOr1zz/U8YsyGbYfE2nbB80mL8V0SCTZ5lewdfoGvCkVji3Lj1ozsSfZVLey2tlZXiAYn
Vi9j0EL1RN+1ZLrQ9USQPbUqBAdOtnTryVKaxw98IgEBgeGjzFRBQ4xwWBzuNpZ/JORjbvfFO3nQ
1yjPTD2YJmnAVtcNGqNMrk1WnhaCvQqR+pHxjpa7ybNCxWej8M20Z3EWWWX8Cfbi+aH0MKLL7Ip6
9m1wwzWxUajf4PlL1JCzx9yDYw084NJ6bZYG1iX703Nee5CjjGurMjpQqh+Fo4mJALLFiAPVLUuF
U0P741It6fwd0JQPiGROv7lIpcJg2QINYjQPCGWuG/fOiiX/bdlgjg6dQl9KiPDR6E/fbFY4gryz
BVl4a3JL20B9bMmpHx3rZi/ZNxm6C6TP8g72Vo59/xO0EjLMh7q+8t2NI6tN3BvruaJhpqC3Qih8
1xNIAG7NFYwQGO5xwQgkXCNufyHuU5l1EVSCZ9toS117ub/RS+Ekqg/mPpihS45xXvIc8PJ5B97x
1aREM/stU51g+um7CqNjDraVTyPqNEaL9ImkSac9rA3yS0x5yOxPzfy/yIBIAOnIaLy4BdoLL22c
7C13NNqiEq3GCg3kZ8YzJHJYWN0sYUvZqRRaJ2kzdUc9CdzXHIPcMpT7SlseALzcxgAlT8k6NVS3
a4SyW3n/z3qs14GQKv3NmVwA2X4YZ49M5qKzuzzZrpxMKWSKThkyChqFFtkCMFwN7Ty9WzIkxKE/
GRXanSnt2iqxcq6TaPXrbtLW2a8+jqcIBa+qkoI23CpWtZ1GKTNq8oa9pPIAzgyPjnT8Eiutoxi+
9P0gq/RTk1gsG8FrJ/BBRnUGDRp+4NJ2BoVVbA8uuWPVp5X/9zwf5l4W3fkPRY7VPLJpZtuULFJg
NV684Mptc/0TgVCzcyhLTRMV0PLL23JyDlYEvWIE99sNTWrMH3DsdLVFDtgcTP5C81mT6tFgj4Os
g3MITgBTp0yKb5TRBlMdNLW4IJofsj36Xz2HWLouxLGrE60otIC1kTnhk44KEM8oXu6gXG9BYhD+
vWY5opN5YCZG0OD13BpZRswxhdIk94kfNJwlSCnPdyBOgOI6z1kB8O/66Io9uoejCmYi7FEYUeOP
8tXiQl+PhjeAn1sg61uwTTb8Eur1AIq8JHMtpYFOwR4kIaNt2gS4FHQe1A4iIFhsAHvUatV8r1X3
2L5yRmDSV19FrMNEbV3i+SVlHuPY0btLqUR47Uoe6Qvgvj7O2mjZVTP5n9Ongx7jxLCnkpXfoanm
MHx9wehU9qaZ0TdZaXwR2OomUfJFLvLoUywjLn3o32h/R6Vsr5nyj7Q2liML9j26SOZUSHxmEvf5
OEty+2jpyHkp+M7Qae/TAzxBZVSa7gpriac3Xe3hK4lwmkmbjlV4TnMdoIrFoZ8la6VGrMbN4YOh
n3N6FAr8o1BhhazHPkoj6c506KQptxKdwSxP1ddk2aGWkCeeP6y1SKXwa5nVLg73LW6TDDFCtLxY
TlxE89yFtFCsDS+8mpchVcbLd7v7eA+csDmfKWMc7BkOhfl7e79LSA4CteogjHhcbyH4UkAeb29j
mIhWMB6KaXffsqAD+MupFviMQJD8iGKHnwweRK69qOTeSgwDPbazukMgKRkjvXayBOCRI6mb1nED
0gObnFFQ5D3l9cWBlFyVsp18s78+j92rkfOsDID/7PEtiIufXXi0oM/hUXebf7KehcMP1akcXofd
UW2dRKwzx0z4IkqC+DjWY4Omo/OM2+o7DroB9OtJ2J6GjhGp0MrEFP4pAtJZvNb9/EKn1Bo95RMs
y9cskus6joZv9vZTL5rJ+k5qO6FdSBxZgna7By4ndVuSxElygzSxwrLYS04vUiiT+787jNd+0zqm
dQVBB7xXfwOUFY5d7kh9OtK1k0U7S2PsGOjZxkkqk1+Pyqf3n7icUF9b/OeHFqG+WbwQKj/2Ar1E
U5HMFS5cY7kv1mtfloIa2qPFF6k8wSNd3iMv8sVyy/2VC8e67Vb4CVPEPIhnqx87YJCSop0Ss5lZ
iNQgsF/3/c7x1tvxox/CvpyysB5L6aJN4lCstTR3lawa1H3qALiLjwDzzAd3TLdhjCu8jUak33Dc
snATvhwQUCLaqmaQuHcStuNy1gTwH2LSZMq9SHLAoUZtpw/hl2IqFGwNnv5MoxjpyjggKY/Otz9X
P2lWdx+uSdnFj+JjRy/ZVSg89BVg2vyc2S71KcQK0UTStssKMeGCFBKf7UNFDXMp0UQQsztyPAcV
XdGvjNZxjFrsJQG9+DF+lU7DgdFeV6Wvjh2PYmJsBy6wlueE0AJ6zYYvMDDnrONaWpq9HsLu5shK
2S6N+ZjP2FQ/I3DTL2Yl+U8sm5EXIA7tXA3OAiPzuoSqfK45fySCKgI4PwGfTzY8N4Vv84KTG6iE
W/GbHYzaVQRDwgJ39s5b/C1ctmFl7nooUPbZTO1IkEcZos5zQMJo8vbrV5SbiEl2+9KN3srccPlu
vMZ2oANM5YGD050jJytNMrqcxPS2DGg1DxpbAbe6sVl0b8bYZoYsHODcgZCGnnT/JwMt9zYi3ANA
XoSwauLC58YyDVEg0Ie6cdWToVse1EhKtDd8bJp8WI8bkRkHDaMq05spWgZFF2NUiwFMIEnYdDfN
jRWiPnq233W+lxa4mtRpjvP5Dfc+zPeVlcC3WYHJtZTD5rSJtEKFG0hcVfpMj3x8wp59D2ktzTK7
DmMNjZ06kO4cxukcWyPQccN4zrd4FblrMT/S6QwJ70/MHq7nMxVpxEIfwh4pKRdF8MPto3uhQuoZ
GvQRXLM2gx2vlrrSvHA+F9RYRlhpSfeESK/U2WF9QfcOWVklvWkAe/1aK07qMn/lvshYbRyvubxu
fkEJKpWgGsbz3ly134g/REbxHt32q8OWcx7sYVDPrE2GWPXmCEiZnmVJMBD/p3TYXl+ECKl+2j/0
ZF5c6ly3Bzs2GTyTgvziDaxJnDTXRwP8iXLWCk6UXf4+Mt7daVKNSleQx9kgFfldyqVFdNFwkRKb
x0B2ummkr8qirxORpJt0HPr4+NOc1vTaYG9RVnV83WgJW3PaxFrVyia09XlvP4G8CmKcYeGADhPx
YB6hMi6E7SSA2FqMh2NBxwdJFZcTDgkHj7L5UnUp7uyajQabsQDxb2MJTBBLW/oFytbvefVWrO+f
UTgNknZrLZT/Cqwnrk327tQI5tg2JWhc90BUV5fpnH19FFMGDOyP6/tQ3NEaVKYLkhcNEeG8WKYv
jlAI4k7A4sYJgKY/llZPHobQ9qyQZOw6zZ2ke3wsG/6ojKOAQ4TEgjpmEfw50KUZG97Ce0BjmhSz
0end4ChASox9ivXju7haCNChjESMN3ZVVF1A0FlHj0jJ77/9UVuzN2DRGyqMQS/z16c6AOwwc+e4
DJoW7NDnskby+/U0OJmdN8vdjCaogJ6N55Px030n9cjTLUMs/k+vofgtzB2k76vtA6s0Pg+NXzQs
mvZetFVzpCZSslc+HLLJuvSjmRB9aumHFQmJyv/dcSqIQZB9Juof94QR7/fG8R9rQHSvSjf/zolt
oq0GcNrHvfEiMlfjwNa8OtB4fL0H71c51ddEeIZWTZ9GEDP6vdaKIWkXDI13oSop924PenRHxEsh
KkONo+sbxc6UH1VS9PAfC3wuio5MrN0LI0OyIsGO5grqkMYHWPg8C8dM6HZYiH0bFS0fo6zzbUKK
qqbzrbUokxb0BXmBcZdIXhb+mVhuzJKoY5zr7IuFCc0HNdAb0WI0VJX+Xw86tUT2ZPQ4BV3PCXfG
xbhql6TQbLmkmf4Hb3YIo2dKOhNuXI6GpCZ1RPnUqB+xVtQEtcNOq+sN48a/tOTdxaYguD9atWhg
q5XQF6T5nKVlMh5Qa+EjSHdIG78KHxPPiS1TDKR/dYcd4j8BehAzyebTnKv2L1qYYY0pcFEmFgqH
eAUxe/uMy+np2jE6VRx0euHqoaLn//s7eRdpSgq+QChHUFu7RDnQx7rnQmUh6DtclBoHR/OcodgF
Hk6J7oDV/PWABjtxlQySlU3rnkJ276JDsTXQ3FJce3jdfN8FSOAGawuqT6hhiYnThA1in1n+LQ+5
vHs8JtL0EPNB9QJzlFrhF8NAUxT4DZdm38N8mmFM4hL+yTC9xlmUc4mkZQvMd6kWha1kpEl21Y3e
grKjeG5pzBYvUS05tXPMMrudAa/HymnYa+PYPxvWMQLiPSBnWNs4hTgFwixCrQi7Hdxa0SVKXqGW
0hejAVk+vhKGyL/ArRoA03Q9nG20HUXk/Ymfl+rXdfmRCAo2LAEVDkvOEJivON5RG+FQ9a2/Yz/2
Kygn0yaQkl+kDOl/dk+ZZ7wOWh9rmG5htiUXf0AQAW4ruSbPwPiClnaJE3cFQDqbnh6GEsu2c+Jg
Qr9mea4cWTVEt5T6EQb9DuOC/Rs0Biif0Q9AZH/v2qNlL/H3IjVU5AEj4itrvZjkEpkstSy48COs
savpuLbG6uMWhZCRm/4gNc6kxsb99cSufdMFklUGp+1dp0BJmGRg9FIgwPas4DWWAg+na84udLbV
OtLRaXjRaaj+K0Up291SlQ7qcu7qU0SOiGY970EZAkpGYgDEmA7qhKHCLPAgD9/baRMyT3OlLRVy
DCzVN8mOoeAYvFtFemN5kh9qudEmd5VTWV3wj62LLcryizF1XuE4/dBZradtGSPMfcN3zhyM3yiI
cHP6kx6BxiAfbkPbH84e5GQsILIQBovWqoN117yrWqm6yY0Mj/czz0xdQyKWZZYdXGMkZo96mBtv
Q31Rb8tuqjypdoXRyjox10wkPrmZ386PefoYhmIyBCSBVYCEQtoT+NpAwX+BfdyhOqRPKxd5C+mR
1DBofMW95+plra9XWovcDBPHWeAzentAsoLf6r5ng3SkihV9CvnzEHwChhTHzS+XiEaWS2e2mjFf
SzRDgdms4GhMsn+tKc/I91BBHPKy63LLUVBVvp3MFgnYDa3RKrYMMuMOSa5pC9vDrwWmziVTBVS4
Sn97EwVtNWlUf930VYDo8trJfDQoAnWmN1cNsFrw9XZQlH0fLZnw2xoj2SKuCp7BXM2TH0wQml1E
UKD83V8Pb9SL3jM5l4LlC8KNHFIV4HZzm3Q7VvLHORzMJPqK08c9gvODDXRqRrI3cecoUhgpFy70
nw1JYh9ZkSVwZ8ILul2Xw8xvpXQZgUsqkcQMIsZ42LgyzMT94Cyz82H1HmiwMybpcvGNjvz/YYZk
7pMmRuSlk5+moL4qqYugtpflO1SdsrfAIKm2+GXHrxmMopTzxaGA9/x9oJ1SLqx19EGconxm4SZy
fMgrykXoR5dSbqru70wnIH5cjKUplNawV9puL0RCC9jooFW9LTwvClfG2RP89HcE/L36/ZrcvY82
FRUg3tSNzYgL/0la2r9KlfMYguqcSaXJEDahOrUEqy2k5lPDTpXQX3bNyrcY2Kf4p7wi+0zxjebf
zSul30+1T/IZCvM5FfKkUZkbDZqlBXtv50qPCVBpr4lmdCUaJjcm+MLT5QI9GjEsSExVpb5TydiT
QnjPQ1dqnOmYEg4JTHlowmYKaYTytTCPckdCeYGrjgGVQf186Xyf0uAXSgt7yUtCZuxW+9MXWcRS
v9mVXh86ucas8fCzSxhYxGkpIWgE4RDJYrjc0LJTajjfR2NGkGBoe4F0Ky4ecTGx7nVE2CVXrrYv
q2/YMK1lDgr3bjH0s1rNR/gX1c2hz9g98MK4xU2LZwcft4tPsHIsHYz0ZrE8W89oNzoWNhaXldhC
kkPUH2tKncVb/AkSuByjAbGTu+ZMjTHEadK+jG8n4hhmaTSzenanqUnnLOXCnxFtVbdDBk+7a25N
pPXzpgoL/PvnD50407SPMw+866hBTXbyMQG0wwiZhUo4b8+XAFNzyEsPKZ184n1omDdStxEiap9M
Rxwq5sPLcFIyoemuI2mqXsY79qQSZBZkOBrchnpQgCoPZb/nTb4juN3L+d8JABwNVV0RleZQsqrS
Y6n+MjfT2wBWRbwkdHDz7V1eV79m9SExl3UCU212JM1jUU0DB15XIhzYb04ymXJfVvPxoosHd8KS
QVMwgcmeqgucFYfbqGSKvqvJK9Zxe6antpdE/pLJc7aa9uzgIda6YOrP4lcVJlR9fbjW1Kr9yalm
GJ0ij1ZhPfSMCOjicqbLS8HbfWjx0R16ooPmdYDRem1kjsbbyhqvy9zBVGi7FPPtqaRUeQd1WJVK
eyOocnjV2XMC61sKjjEo7QaAVK+gQ768TgEWWRGH4UMg+YXTWgbzJRHq5mIsJG+xH4VaQP7u37dW
53EUEfLqs8zTSq8H85x/KWmfHidwfwseIAkDt1KcQjaB0I1zluwhVm1w43t6ncAGOKME0qNn8Z3o
5to9a6ONsoi2Mg8toFvntHQqjOCpqmf44sWO9hEDakzGpZEpE/Ljbra0p+oQYQJVDL0c+ysq++7I
PgYndfD0P6DN3LdZ0IEsFWwC3GnVR64c9ZjzhaKFFgQyPEXt5d+VK1+Af2rB2TLvQzMhQJ1Thyqu
WjVXoYBWPPockH+dYJLVlUjeerGSJb9whMHcNe2pGoJrca297o3tS6xJNoIvdTN7FCCh/8tbghKu
jyOfeNtHHO5ADQpQZ+roHEcCZpFzdO3nJ7zZqTuN3YeoZlkXvcOn+bsx8T4Dc+WZCpiVIij8Fxdv
fgJsuCL+rE2gC1laOoHrezd463jqfCkR8iErtRv6U+gVMS0wtHcJ2n8QCMBzOXkn6OwXHBJvANUg
C01au7a8rimbV4P7Gb80tqbwJMeAF/00/3lEs/OLL73PRmOdIlbM0fYXWBG2KHsaGwFVR7HXcRSj
oUCcO6TsKEnu0zL7XZzynIN4fybLDvCZ2+lNRS7Uoo0+PDYqLoF/qqEIjjy98eCmfdEyudZqPE2g
G1VQFACovi+T90KFSEb1UCNSzJAQwtwf7FMSUs7N3THN/0XvUL7SJz9+qjIi5gD0IJBzfgUfxZc6
1/GRft3phvOejzXpOPnEuWI9Cj5C9tjgTpovpzqiscvhrTqDXImQxxv7RUg0E0l6gNjSGaMf8cQ7
2oyKucimpf36JzxS5hq6r23gCT/lIe9qPuRhQZmRVfLy+KR9zZS6m+11exZzuguN4eeKCz7iBlgx
4rHKQGJZqMqe+rPo8PczfNFXW1trk0/sW4uepX+xkC/ILBWA9mhGs4X/PYH6Z3fUctgH3/IaXOkg
qbAl1sQNuJPS2YWeuHIC/YWzBTFRuoGpXLCZlDJE654MuStSxIF8BpWrniAW5pHZNmELwftOqDXa
im7aGYOEIv08gWqgC3D1AUjK91hktgUPI0HVqfolA4QgK+B/aDBs9SVg5lDLtjO/2uB6w9j9SEWw
CUEx9PpzVHhB/j5PdUqkXahgCRCAok7b7mz+Nt/sJ/w63GKXAISj+4cIcmwjbYRy8gZ4PnFL7myb
ERJCzTNl44Y6Y2lIwnOfKh9WlJ6e3V//7vg2EzBDjQ6UOfId9f2MrsoSiowcVGLLOQEe6oS8lC/k
4ZZXFfnrnLotN5XYHtCV0scJieRcm+Ln9CPARYIXsxTvDIGwKcIGsOUsmfFAVsF0gicNax4uzWpB
koCupCkTE28pLESlFWHH3J35urUZBWOcZW1kPRSuGSuwilF+J/PqpX4FpAecfw8cyNA6WzjekYma
u5oXgC8yvGiQSE3h0T9SyrVgXFpoGulBBUd4K4Ce77JRPBLktG8Dfz/+wZCxRSIPIPVbPNXTWnbv
Ek3hhguK6JN9KlY91VamF9HdsiSTcfZP5sYQ9zZQ5XgrF9Yh8Y5zIZUzpr05UbdycmxlV3syV5qp
/aMUuPcHLUo/+PueBuS0dk8v3KzrH3lDWjAaEBI7tS1i/aDC2YkFWPwAueYD4sd6Opc/Zr25sK2T
8yLvnhr79CFOWJDY0VziQ219eq8R+X51N/BjycKY8/aKPEhI9L9U6xzX7JGXMxQox+h+1xgSZ0n6
NfEFC8CtRiYZhDA1QZV466jO5tdpNdLfXMniFY2HlFjFQ0fcRDWmx3R+UwYyob3yWp0LIHbS3Zx1
ZXFSZQ6x7/rX5RnwcFhtAvbV8fvmLmSYjkVI6rWES+rjKF+Q9hsgL4DMy9JnWNKSv7FI48D6bSr6
Lym4Ac+/EIZVlZ9EBbcNDduROj92gc+HHf9z16lgZZ9qC4Ca1kBFU5AvDxMEFYe4uROZneHpemBE
yf5tbiTMbNZWUKqRJjtp5ruiQZEkrXu5bjre1YS1a80buk55NShieOfbx/ZhSbj2J/LK9VYpEubX
6DFLGTTmt6s8KsHPc/4KdR73PvumAcIXrypSMOSNLPjg/pJ7sDwQ2eICTl8Q1hwfqqToWg95Fdqy
Q91cEyRQdibSP747Fnn0XpBGUC4gTv7Q1Az/QmutCGxPwlFoTCcEOGCzVSH/joV9EMDxcXgv71ck
3jmMYA5ScgnUJtqcAFW3Lk8d6UT4OlZuamlBdf6qEwDo8OyzD7Jf7A43fNwpOq68OEMvxytjsAGX
Kya+bd1DmUoOrkiTOIF9CyuOJxZ06hBgfcJQYf0U5BtnCUm+e7yQUoYLQ5APVwZVHBQ0r2syu+69
FeO/EB7Q/OVdLRrAfpBVlvMXIDKzXE5Zdugsjznd7qE7ctNdc687y+yEN+4unKn9ZgHsekLuIsJQ
5Hkdxh5TUa0m0FzytFVRzVz5hN+9Um5d/ocVfw2SB3IAOTlJpZTaoCwuUlXl6DUZcunEJP6fWqyl
VV4xNwhu+X04PSNZZ2TfDEQkili05cqr1sY0vtF581UdF3CyNa4YjLcugPaChj1GR5cQQR3FrFSD
T4PTvdxAaSyOEcXStRneKYJcSAB/qIvsCADBBx++4cmEon0VDAg/Oi3aPAvcdmM9+pGGh/d0owfv
pwgiGgYX3LIZAX/SEsh/HkEq5XbAhO2f9B634aoH0e/cS1G+s3JQP9HGufsIVSPeD0UP+oIDH5vz
MziOSncwabXLgWbYEi3S+tARwzhQt4krFAwJwCw3VOuEQRS6v1SOAm8SiNvlDf6oFaCOC1F3ep+I
zK1soJEkEtgwfJFqxIeRevJRW/beJY50Rysi+2QxhNJ+2Q/WNwQ9k61U8DkN4/2F11SQFFy3E5E/
hjuWyxCODOUgMt8aHm5krPfailT1Gw6HjOXnpga+qFO/h8Hk9ZcvYhN97nh2jVFhOIvSQUaKycLr
NHWLXohgl8crE7+c+DAs9qWa0oO/GBvG24YfnU2UY8EsuLkKlQBOLsGI0AAJOSnlTQZd7uNiGzry
dpgEI5sS6QHTY9kh/+uK84eTyLPAw1iNs69XQejyKJY7H2nOkL6/nNj1mOCt1hoZJ5QLoSljjgHz
YAvICAdm76t2vff0x6MYKkLfBaw109MnWB8F8EdTqKkJ9XQ4pDDJHHsqHn8uKyy4AMBOV4awRqkG
dcanRH1c5W6jDX6BWg2poFonTg9Dgnn+NZbZdvfEGBXZVBH+91mq1Plwpk9VRgDJ5lH17G4joZOw
nySzczS7TglrXTk/pmu8AytC55ECT0SfIYKf0AkjQ+w2jBA8tZVq/T7u+Ml1nDESmZhvkYurUvPu
qk3zuCbbRBdzFPbTzVB+HsplnJU1t2VNegqNekyk4Tn8pnyaMcNguy813kxxxbk8F0+UjkIZdw3B
Hn7h+Das2QzES1ZQob0g2dB36Tt1TqlggVbyiKGzau0TIygqcogw3Kv1WUQ38+CUnFOsFuIe0ifi
mFnMEE5rvhLzQ70qhpgJSGzw0fOdVfP13YA155Yaao7bn/e++t6X4j+nJ5q7OtJcIkdg/oNGj4av
7zyUncIezfbp0uKVDBx5knYBr+sP2XuIxAZGoK3Hts+5A/Oahvw9GfBxXAaZI5B1gDwjJ/4sDMpv
CGv3L4tyrOyN3n1AUK+CrpIj0BY6MNt4NuqqUYtscTFmsB1Z9znAKn/3ZefKoK4gse0H2Zxdx4HE
1cglsep0EY1kZI12L2OoH+N85YcG3mgn3fr6fW7AX21sI4SDlcwOM5/hP+oSPKvc+hdIgeNu7EFr
Rqm0pOjpNgJilmgEORpSMvJGFeqwiRd12f795GhoKo+TF7Jj4WfPMJFBJCsPF/j+aRFCjLhDG8Ih
ZZKpVKfuac0P8bKdtDRwuCKzv8105A0+qwPrwmLM4kGzU8TVQ9KxAAtNZ5rQ+2OUB9Nrc7S1YPmY
pbcdGd6jwVLSoGfnlml+vkzM6by0STOS0XmgmxNNlgIMaHOlxr++HnDBsSKlYd8mJwj2yp4gcG8D
dEO1EDbok7VW9X90t6l15qb7lWHjdVlm9LPTdzwB14WI2x6azSDzfpmEtEIU6U+3r76OyC1ZHgMe
fQLRdTU3g4eaIPOELZktaTyU0XmTPFFdv6Yx03JZq0lW98uYa8E2WegR/O1yB6e9dDUBdF3p16PD
uEbZUZNpMm5xaCe2CWr8c9IV7SPMU3YNtphDwokGo1SiRodzYql+nRda+BdDDnLRhgG1p+nnG9lW
GdVSkXLVpd/2kwpL8bCZBc9KAphrWne71bSSxbuLcCxL4sJGNigo8pPrUrTaUZP1VH5LHkM22WHD
iVNBiPSEixF1D8zXig8kO6ZxbFhJFN/Z87EwU1UBHbYrX8hPlUHVgty/lk2JI0/Fq4O3eCgx6f9Z
1ALbD20vzXuTPaEeOunL4mk4Dz943GGSjOTM4dM/fISRfbYsUBILMCuTjfT2W8YcK4Q2d6GWFwFO
pN2RGCMHC3BAkdBAdEubEZ8GiGVOceHM2BexL2uDAZEMeCBRh5VBX1LH7p24xHvWrbdtTvlLFvyp
RbOl6fZi+AgnuTveyGk08ovO3ak3CnxM2ynn672Jn6WPJo/F
`protect end_protected
