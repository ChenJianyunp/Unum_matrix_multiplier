`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JcMz5zej9a1ZiWy011/KrbSm5eLPKKzlxyICi2hv0Xw1NoSTAO/eZJwAuNjKoogKS48O2dtJwuxO
WdRxk2iW0Oog7m7K1TYSBSYhELLcV/T0EwC2D6xq5vetURgTYJm64QyRDiZFAEQMh30iGn5gryBa
BfpuRx7nzG8pgWXfIERJxS8lw5UX4flVF0P7n7OW1G9Y+gfEHClbyJCZ+PFe7cu62eH/8raGbiAI
onroh9H76nGe2kGCOldYBfRkLBBv1lrc0pTM02hDbBAMBcHUSIKozLFkzS3Do9zYCB1C/EDjiUDr
lDDEILyXmwFB2Qj7GgnGIgXDuMe4p2/UdLsamg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 111056)
`protect data_block
Vj7fykTb2u6mk7Uldj2vYJKynKw3evH49lWSzZEX+2Wpj/hXgXkHXsWK34C9MOA7mid9K0vI0v/9
1Xqc2vAPBQsC/GY/OM/NxKG/+KJD5X/7ijwV7d6kR6PDBPYXiFqjzM6buWfWSENdGr4ZKl1LqO2V
AhL2djNHLw8rDtlB+yDTyErxeFaDqqeQgXb7ua2Cj9E8XF4AM3t6BlL6XpCt0imvIfNshZyzSb4T
ScZQbdRJMhPjgt9pB+ob5krkWpXo57Eby7UYUfPq5ixOEhHc3pKrvVihOz/desjXJHUntWw1zG8Z
4G0pyUqbR9m0L2YRBOHC1Qm1R/7wK6GEURcP0s/h4D1cPCEeQnTRMeIt1X/pRW9bJQc7AUP6Rvib
vui9DEql5cYeu17ApHwy7sVV+tsN9Yv4nHMnFWyDE9qeb9ThWUTF7wB/LOrNUlprX3U5zIehsjXq
OPclTNdMxQDOUd8SP1ePsAOsIwV8RbdNqJBcGoltYLiuIC+pCB3uwH0lvRNF19MLBenizMQZDQtc
N9f6b+DQVDZFu3HpbgOEbxAFwSd2EFfsmLYrG3NdC9apJYBbBKIT/m1uVH3NE/Cabv5WQEv7V+pl
DLso/E8jQo3KeCw5Co+rr/3A45dP1ZHc1pILC0yId7GnmhoaXZtKUhZcdkpCryaEqs/z7y6uM40b
J8NiF45+rkuLHhC1pyMEcnhR1z5U2OUEtMwwIMpnMXiv2+OYJtuPp0TyCVj7EXAyqDANh+/Dkkar
VbKceTF1z+FVC+SWhT62CVNd8rXMpAnEna69olR4oTvrvbrECqMJGascK5bJe6svh6YnqRXBKvIP
sAbyXn1EyG/pL4zCndaakpNF7SoQfS+hqUEfElfEhUa+f0OjiaFJ7gEoeJi9lmqkl+F5c3oNofSN
XC04uodRTskAIJcqOH556ZEsoka+Jn3sOwVRAlRvopVF4yolu5kdlzdb0nI7kSPbz1040NbbheAt
FfTIbGJ5cP/c4sIrhH6/e5DVo5PI8R/ov3+UPPLWjIVTNIDPR19eyg8uoKxtI18kM9eHIRU/waiH
pFZUuWSR0P+tHjR1XuLyskXviFp6pWVCnQGwrnPaxq61ckqLjhpQIeLbRLhmzIrHF/PHEo8+B0Gh
xZQ2NkBOSnV5oUy/b7MoYmG9wMDO3KghE1+bZwan+GDxC8YCNDLtmh4Yu0Gb7acmngNaBf/7L9py
lsULuEU2unwNVSYbcIZ11wz/5d8ekCJJ6yE8rSmfTCjRV5wi/LCqzXUEUJRI4UJsyievR8cWhHcU
iJ0ctzTMEYfpwZlcaJHeOHyzGowAOzSjYHp0Xa5u0PS0XHa7ttP5rXLovM96PJdTQ6Yt7qB9AQv4
MmnwVkB39aGbmkzumqcifYcwASBtXnuuv7OjvFmJLWKKYR3MbwU0m2x+sDSpCxGBTBVmNcgrQucf
6kjUvd+p7PupT5dqJbC092anus4c7radjWbzO/q5It96p2HGznUZCKwqeGxkroG278XnL3umiKBa
Pung50Tsp55ohBTL1oP1fWmufgyIhyM865s8+0d4PLk3VXKZAI2C1itv2Nk35EcxYLbVrksj4e7j
0MLPQlYQz29pnsVjLLWWiqxa9NuqsxKOk3HgBW1Kan/ZGxxxQhuWMUGI/+nWO1wMAv/5ryYifLo/
jx3PzopsXLMn7P826z+RsfiL2C5MBj6wwcsg9oCgJuBhKE/YQtxSJTI4QF9SILC3nkyKUkOLG99R
3lLA1fU9mHkpXINJnsPnAJjaG/rSfACs2h4plzlZ7A03i7d0cmIXoFsoDu/5D0N8mvXoi+pCnM2o
Hib/mLfSlKCK/cwHRNxCp4zIHqRZ2LaGG4svKWvYa4KhJb5jwjQJZBesv9D5Mjihj0HZP1x84COB
c1HiE42k0JgPIb7D6HSgI+Y1Ks5ZsJJohRMJ88U3wYnoOh9LJMUFTUfHsVQKJjFN4Rumc/01fPvz
IjQ+Szo8PBHGFdGJhZEF0DgB1pi4ha7iHd9NS+22D+quvt0vGPGcBdlt130551lDgiqWfJteUGWx
DpUb4XdkNSr1JW1b29GmDxXc6bXRSRN0MFPgxBBZTOlZEjvnIBfix5R170E+LBgLGVyP7G+FlKwY
FoQnLSsltz/owPUNqY+FRWLbPPqXKofYsdatDprycJX+wPrDV36xbqEIPVwKFD37iP0nU/2hxSjV
jRFVeL4ncUNj8JKT4tlQN2yhK1jU7PhRSvIlod1U7UhOGdiOskrIigBvLdzmSbxv+2+qDan+8BIe
OaaBQhjPbpHfhQxvxFOZadzpNrG1WEkR5Uf1f9vwKA7bRFCmfJHHKaB+kPfmFvSPkvz6kQBZm+0L
kqGSpgQ1YyStqvo12dR/lbmv56GJRElOVRc81A7yP7MqgbvLnQWtxJytEO6XBuCYnEC/undguN4C
NiKtnwqFVFH9EDNZTdhb8WAJGjwZSJV3n0hIweCN00XS+7njKcqdXSSdGn68LVgBlsC9KWX9IAKt
7VjqkI8CtxfB3lTuFwAIRz6Lf+rMj7DgrYrQDlvYYeQ37QPPHkzR3uG7U2BR8+ai08NnTOhnEA1r
Ngp4YOmnOSVZfOaASMBSU1c6tG+HPVfImG036v/wVsJA0CeqRzp7xYs/EGpE+xDOZrMvEcJfzaSF
wzkuMXgtOp0aecXoX8SWw4vhqVXjl11tzZ1RKBJFJIc/S2DRuX1RmahKDbGRgCAn3ehYOo1vy2I4
IGWmXJaVXHmqdRJ7r2sk/pKuW+WcHDqmH2glwCQZTaLWGrki/8Gv2cmG5WKNdjYA2js4DWXa9dCU
slvGbRDmHFA/YCzTr9kWp1xx+0oHGhO0Drrs/t/4+54GApUO7eML6PwNR1649xrOTDTNTvnB9K1m
ScZOMNRk/+BnyYzg5QjS+mK4rnPz+DJ1WOGwgANJv4YpgrG+YYZdRrWEpk1F/kyJRkcCd73IASbY
D+fUiH8OedXdEOVgM/9zplG/Kt68RG2n5oXZG6g58FokI92pt1Hv1EBh17LYAU2LGY5xICWv3z9U
bd7jKsn+A5q7paJPvuwoOJ+WUzVVodGkcEamxu2anq+hVOvuviyMRHBCuNREorbR8ls3pS8pFnUe
SVd9LojdiFRgnMV9S/nhJIzixgUWlEqiwQiHiiNNAg8Fmh1zWJHVG7nGNM6pur9SAT78WzTei5o5
uysdTHZj5bRS+ntQe1h82qjhM8UCPT4AL4uuMZQVWX47+FWFQPKsyFpvKxMPB/okstmnlWBsyZgs
CcOdDkEkYlpK9piXH8H9q8eA2fpyUiW/PItzYY/YpiF6sxpWleft+tCOZyTn580B9QOyk512opIn
ascakShIcN78pDTEsVzTwAMnVX7sqaNLLrI67CQITJZy8oTfITilEzqKPqMnxaRNMbld3QgVbF7T
R2MbGdNI+EkTZuKE09qN4Q19SSBWnG9iCvU6U07WilgvfOctAFetX1afw6kcs0UKwbAngm9ZEE0k
5zKQekyzXd0FVYpbfkzx+8PcK0N53GOde/iKecGmAOmGoBjXmVTAunEnSALCqIajsUReDTAH7ueI
1x4ufx6Uhl1y+7WcF9e7SkaQJACRzQ0jyt3n2Chj+IdbFx/C1d3HsoUOB41lEf7R3ho68UwPvF3I
2xW7Gx9MGvnhVFx/D5nze+ltHVbRBQy1Aji6OABWh/9jPWE3L/ljQoz2aQxiT2FkINczxzCykbnp
+HQ9Ws5IO1chUxjL4kJFxM0RpRR0AvqQdOin0LIGRy+r0+VwGoR8vPsfL8BNv+QkPOaELD+yutAb
8YTvq3/1lKcGKkguS9wjANJ6qDcHn7AOBNPA0KVrMYamu0rDn0+Sqg05JlNIlH8cYXeE8bRD13Yt
QrgByIWpb7xxywkgEtfkKrO2oU8kTzyISbEbyBquMOBqeoPyIYLyfkDbFslV/DX+0vZV5w57F2tB
VEHclkareMCKu/Cq6n4YQHW7wU61lzkgIHA5uu312BIhNbreReGzFh0JCj4TkWFMXY2xf84kX8Ok
pq3HKogx6rPWvy0AtVo/bCexrSBP5ipY2WhCAn8OZNSQzZXTlLYm6nNvLSg3uj044O2ZgPHllUSW
FJtdIn+GoBfarDZQnDKPsEsYSkD+ShmPDXYhijBTvG3z5wLZZBNmMHqeYTzeudDlcDrLTQ8W3N1Q
8y4p9L70CBrhsHhqpTHHq6sdIst1hb4cKRyClIJ+EOt8HCuLWcIVikXvbn9UxJy/Gegm/fiWsX3w
AjiQpe+aDgUTLrHN6f8M37+7zyTR3Vru/1omhHj+gWe55wPFZMqOXnKPFiX6EmCdVBZQ19ND34P8
Z3qXw+1T0iM96WRqRr2/Uwo52jDlPqZOPveCXr///bL9HzqBjARFpwjmkDJWVhM5ENWLLHBijxaU
yjYsVjvhlspN+999f0vpHG7VPrPkWMRW7V+nnQy0r8irUsbZHlDCVoRwRl7N1PU8Nc0B7Mhtuqnk
Y8iZLF+w3cYHB6N5TviAPj/3tya08z2mxScidcp50gqFHBqCV5pkAHo60BhbN4KnoBVy2eBhV/us
NsVN/v8PHFNMxaucY9aVnnyY8KhuZ5C+wJcwbENr93uYcnLXPsdlHMx5YF54XKpgWAeL5+UmMoFr
Y/ZbSt5WMXMEdtSmBms/YdqzjxUGUiDIdf9YuVfoVgIB5ttI7U/w016ZCVGvZ2vsGR2VZZ8jg0JH
NNJ1BUtIDxLU9Pp18YC5xDfxe1AxVcISNPq97Ipl8s4ivDcWVtLcY0MY2horGWmCQQQP3TCNiyot
JZgNJ86IWwhA8OPP6lYu2lhlwCg8q31EsrTK7F0X4oC32/IRYm7NsweXn6Y4oj9m+J/7J4w/oHbm
eSHK32JDlKxMSO/pot1SLSBjNoq0IxhjyalW2shHNugRjy8Bpi3qqU52GcO6NX1pMTL77SUT2Etj
YVkf3X09Dv7PpR0X9+qofRnN/gWrx3zJ4tH56nKwEtCdtIUUWg64zDGkX9GaNoxgBrNBgW3XU97d
khfQrDcKrdLYVN1uLMN4ZxoFC1J95Kh+cv+ifCNXpzwO0A4bwaYI04lFDyatxYmMOg4f7CiCFjN7
8dlV5klpXrSW73ey1mG5YjzFMFY/pwCaqi6qevNNT9+VwDB6glWyjnQbiLzHoKb/jBzqooHZQg97
wKLCifWAAAK8+sD3wd6XIuNmsR9FryHifVQ6kzImP5t/mL6u+cr3nugz9L3SiUTEBKDx/ndUF5W4
2knDdGb/N4CjGnyYXG3lZID55qt85lLSsir25WKnU0331S+JmZCqzl8Fy1d236kNVmSQlHfo7Zw/
X1v2TEytUAOh9p1NMN8fxtCANGXibYSlIyg+1DOkJ0oZ6nkmbCX+X8KiUCuoscm0QOziLFYY/pE4
va4o4RUnsM7pNEgzDZ2RvRa/WmiHE+YYErvz5zNV8DvGotn1qlOrU/FMiW/RnSArVaPu85/BSM3v
r4liQyJ1aZBVAozm6zrHaWabjzuv1lHQngdK1Fhz0ywQnYokgFyWRYptB1VtcoNQF9iYyIrhuSgb
OeWULCEbtHpbAMafZnI9jtL6TOqV6YdoBZIRluK57CrjQhr15PXwzlLzaPfMthVCvRQ8Kgtml2kE
Obfx6ynzrhvsYLyErpJl0TLL+02BJxlm6BHh0FFu2Ma+fRZqiGcq678gW51leDECSdPxvXk8t9yP
92d9ljsc2JRGCG9g4zbuEqQHMeD71B2WLY8FUqrb6ynoFjCRK1OpUGGHf5bpqHwIksFUDlcu+0tf
x+eyAQoUFDzndrKXWZFQH8Njic+ytZrIVilJJ/aj9E6oAHgIfa2lrqJYIsswxyBwMCRDheFi7wol
EOchgptWIlrrtliQUt+zTfoqY949bsBRlsCtmNnbxefYBVknEiSO+C7SO7BrEQWZ740NEBo0PIJe
jRi7ZabZYSQ72r5F/aBsV1U4xHG3s+MMO1F0PKm0f4T1MZaW8EWpEIs+n9h3lZtj+/4qpbT+2OhU
potOTR4ux5DPFS2RbuxDV4Ho9ZB/qVSiooi3gXMgInha8HAOzG8s6781ni8LV7aeCq1g4pBumtNn
GwKxZG2UIeQ69t/6rDSB/5jXJRA3Kl/KeE32KMj0ojjoM3j2yNL7Pboh8hb1HFgYic7kVvsigLxu
sx7/3KyhO0j1qhPqCkE6XKaiMwho+4Fp1f0HKBhOt1XngbNpjmTAETEV4cg8RV2/kUOlAWFVKLuM
hqBsXNqF/XvbtgzI8nayh/nxWfaSW/Q/+aF+OdsSRAO4eU87mrjcZvm7qlJQva4hDemIUWlQ2osA
Cd1HqzUtNoUCtt0AooNUdQWkbZKuvdbudvhDh0LnEn2hD5AIXMh3BXxFQkoFOYoOU9V8GGfDxPh6
/zxidadT//VcInmDiMKTn2uOC61RaR2T5jBm+4ahxDzBvbkk81zHQlIwlk7/QFZzxrxN0IdJarAq
Y3jtGSmqNpmrfBzSdClrzRgZW4YkGgaRHsI83kW6kkCQZ2WI1UqYw5kPI6nusulfsXHthSmG/hsT
rV6p7PIMNmN7t9daBa/V6dG75Mabb74rUOmMrpWjXWH9PEZzP6b9th3muD39ztks28wqXM0t89wK
U4ctiUEvnNuj6ZAoPNPT2+9jlx8BS8ecpVHwfU4srwft/8ayBcoLjvxsVb9cFTQPTdjyNJWcvJD5
ZipYOunZzrVy09JLK2XZ/xDHcgcDC1sy9QF64kDDQOnw8gqoK/nCZxnO4GUK0+5MknpmKR9rkd1b
sAK+Lc6qe5zLgggB4CJQL57HOiYDDeWkjPSrtsx++7rf9SHe2Ug/nspGbYRaaJdKZhXoZBSJunFo
1GvikYfYVXXhs0rIN59vxXdeVzE65hU2lyIxJhaskk/tmjhUYcqj2c0nLcyNpH1tQx37pm80PWOg
9wcKDaapJyBoJ6N8+zWsNDPO6R7ov23uk0TGDCatXDMfNaXO4WXf8FTMLFESnXiN9IeQSfs0fi9t
CShD2KMsDTRiI3l7kUy01NLs3CnijRcCw8eUVAejT2BtNj02zdBCfDWEYowJ8t8Uqv+ETcp3iSYA
znAnRh5fCngx0/zYh23e0jDfBX0WQv77RTHEyA4aWk1tNn/77S8hvbswB0TnRdke+uaMimWfFdum
qhhVt7leJXBKp8w7P3B1bD/TE9HsyzLrdbmRSi6HFPULmeBhlW4zy+N5hVTT/oPP1phbIkO5+nWH
f3+YUVz8+lH6cVPPNiKShjocPu3QlalEUKZ+in7dEjuUJMK+8NDOQVH1hB4IsSFDioq2YY10u2SP
pE/eU4EZ9stkH7ytXcaCWbA+yWFgcB75e3Tla/h6ii9jJQNwkYMlF+UAe4qVX67FyuKw8ZuKcKtA
2xvUyIj1lCQaCZfxMeVtKQZhaFXaZQ5mWd1p6cLkXZPwh4yOmTzhQMBGtMTXOn/BUrS983Y6Zmpr
exZhxTTTiDlkNdglc6qET82NQPjJixNDqVpG5Vlhw4DQswevShrgaGIJvwbJMbAOahWM+HLW0Aja
aMAjyIXwCXDDi5KNAK+liKTF3kqmOq8VLEOh86rqDIFqz4+Qu7eSDuI8PtWFYVcarmbfbiI+fbZy
p8v5lYATulwcaG8b+SaSDhMJs0YHfuvBYYHn+R7ZP9BeC/7O0qqrsBJ3DxiJpE9dhGEI7fJJDE7a
Ed1ytrZ5fBM0VyK1UhB2TYOXCmeVBe2dB4lL75DgD6oFLNCcO14RERhaEkbO2IAWCNVdBo3VJR7j
tTjiUoH9WX4DHnYqf2EZCPOPkIgcDosQLww5KyZtrHkUs9Lyw5lKPwkZnxXzEHMjt+fdSwtPbvm1
sRXaiAC8P8o6hnzbeNKvisnmIspPQapEL0TDG+348r6bcQaXnw3vNyk23v0rsmxhupItD3hZbfyW
pC1rIZVijF+ba6KodYPMDYVet8rv78v8rHRp+bpUD++qoSY+tcVpWb7YqFXH/OWkh9+DMvYV67KI
WgvSNFIS60sQPNCUrJuGjZiDIJ7/Wb7tLXr2pQVvYfQb2x5mOZi6NX/S6nI8L7y5kw9zbrNP6CvR
aZarmGNfjLrGCMM0bA9lkRXPTdosTOANIS40CU6mKCSYLE9v0fzT5CRfD1pPWHxcdMqTpfUDg9sc
dILe/PNxAzKO5svcMQSaHZbiJMiOVF2I38AwNFPhyesK065gcFwf6LZjnnIxthd8gfXb1bmLtxz8
sUzb8A9Lxm2+Ts8+HBZM4aYBTHKEGxcV+GPMIrfilRl3kp0PPZUOQajdoT+9S+BGNcohcP1+x3Cm
bDNBXK2btKY5hmFSvNn88IbRwqmSkS/W6LCPiBRJM5/is9DXKIVS8lVfyzAHjMKalK7NLU+F2h7H
0fbkppJKEQbeQag0nq8cIfpzvTqG1vp0qkyJAbUuRzp46cK7PzBgrRXNYFdh7hMTt2yEAanQncPt
R/GsDgeR7DF+INY2KXDzUl57iwdF6O2eY6aLMMLKmIIeKCOzlmlbH0czf4n0M1t0HtdrpCm578R8
/a1Xq8OWJYL+6WOhiKmuvvfZOOQoKElNbMy/wmOX2D4e7KXlwe27hsPKB/mVxdtY3VoHErmo6ZnY
qyI8mJRffSjVRhdBd0SzMuB518tm3StlQS3ZUjJU3POYb3Og8e23VXybY1KKvluBGqW2aetCnkio
+NpHMfmDL5Nl2pwo1NVornwy+owU+qmygIQjrR3EbRXyMw4/dNzORWOuWlYU+aZGlM5Y/Yxy7FqX
zYeKriMmaLJJRIvgRH0FrzK8UZOQ2Nz1kDgwYSI/XnJzTtZtlYEEJK84/9XsT5sSpxgORA4JY5oq
IO4Im4RJcSF+4e8Hx2wXlQcEdJinVx1OKMyspmNudNzLBag912ZHd7WfiCpUA4FsOi9o4/aaw1Y2
UVnu7J1qsECbhRRuMhVI9hqhWFaE87wdW2u0X4S/kh7YaEc8h9jV4DOFdQQbpuCsulcA7UIxw0w3
Kyl24q1xCDexCi/5hht4JyAIhILdp/hqEYBi63t3QNGyOlKud4/MVXudm92tCd8oHUzzwUff6JeM
96i6RerwiCcrNIWpxP39/dxuNuJA38bOR5WjGOVniC73LqBF9AoUQbfe2USWuge83MOwAxi2azvM
1NBcV1H7YWF7VhLuN7bFnIWmeczd/I7N/A9aOQT2ZjA4DiN0RJaRB+pqr68sijKdqoUAZM7JfFJn
E9/fApiFCLurXXPZvLXh4jQxlum2GJY4ZN6q2lwkmFXk45FjnBkNrktN+h5jkWlJPtfNJotKZpaX
uREPC9fYM6tmKovKkwkjkzfKcc7xIOpM23FROnyTePiB3dA8dEPDzhgmwXA8TivQpylcl7i0jMg/
N8ewkBlq2z3qqwsAvbdYshdaEn/oP64lKPQOvnUvfP9blpmZL5+gLLO+Wp+XsyLi+N4goM189Bt3
WftCdRkG/2ATr2qPevlALIzjoFQK+dZxg7TN9kG3HkOBrS5jDaWl8Hddt9CGsKo2KVtsDsHe0bGM
KpSs+7CzjAf/J8RV0d9KU8gd3OLLiWlp0w5bizvQ6P9DIEKShG2T3LMKx3HKnfm04FSWeAtrCahs
/BqyDjVqqF8jedCRwhXY2o8b3zQk1isYj0F8chMTPw1za3zLwi4YWIv4puO2EYeBTL9eyPPR7mTd
WLqEVX5Jf7DLQ9xFG7TfftqEGQkzRVnmnvAxBibfnFMXKDdh/MGEpu8PcRqv3BZE3/+HSFhd5OJH
3pcfK85TtfVzsUd3msSGqHxPoreCax15LP3/opNpF6PU7ZO7CfbagXZmbGklMlXe+oudGGw2uSBd
qwQbyA+faKQa3voLP+kWWG+VSQegJRrlf7Ehj60NDvYT8Va+f+23JGeMwJRHuODvZqdAWWI+Sgdz
dT1E3JpXDKLPwmyyFJt6OzR8V7/+o+DSFUcqhj7hvNY3K/bDNxQsrV4KvqRheuIkeuMOFH8KpDkE
jESAG6gQnyf+3ZT78EI2NKsmgKmRJVysN6tg2oeubL11QL6SW0nRgfEXk794NPLvFjASU3nMbGB2
K3B80qVM2lxYgSUOSTk2rf17usYk8J0UZ0vFCjdIYd5uX9jO/5EyQdTDWrgvVvUNber/ncyOMGCR
Pma1AWsbs3kp1IiDN83RgcUKSt7RQGCKCfqnu/t79h4nuUUcCTTtbAgkH5AidmeLRGSv1F2251sI
qpZW1KT2cDMdzSchx017L/tJeMoG5MyfyofdAgsASdQdSnU/kzzocvyP8Yw1KBBm6WLKV3YBYpTv
9iJCF0QM0es8h8wB58AxDPe//n98rSt/naAbT93WjjpTIk2wW8L0j2ED08vk3vXLai+5LY018m7t
IsOuwbMQ3EhKuzCeIcQ3GbQhfpDrCG0XxbSfYEo8EQvk/RVRMBZt7MwuTk1W92Axa91HxP8IRDcf
0oOU8spGyptmas7gh+Yea1k3eLTg04kViBrIrAm9GdFUReivO7396IrT/b9MzZxK3mWCR2EbTuLu
39fTbZIbbESojoWDYUHbZgkdbPrbySRCatmEQn6rIi59z9hsHNJ1LyJvYr99C1kRfjTlwcOMiDxT
FZ6ofV4mASYQ2g78E87sKMWw4CVnnfpZcLaiNiVgQ4Atvq8XVbSWpepLU2R7whffYipfBoWv2d8Y
B3a1L99q2smJ/zJBvzh9yECBGvEIbq7DN4VAXe/QsLfJmTaDu49Lg1mwRr9cwakGvuYSQqDVBQgL
9McPX8enWKP3Hw08QEsa4JdWtRfY87D1VW54lOPSknq+Hfumnjkj84QpdCvVcI+bFm6uKCyymnsM
eqpGpnIJnT/6j3Z0k1slrV03GQ+Q0HfFsSJE3+q5NHYBc9oHXP0BTgkZIJXSFIcfs8tFSim3TlSg
QsAonRw4mvvwfUjvte9zQVQQm3hQnMt0JU402ZK7JRHCR3N4PznDyVuT+j1LUFBXYT433pjtK+WH
U0XwmsjEDDzseiA0qbPXHNZVKNIJZIzHoZC/gh7XJZQEPazRsp0yxiI2PC/serkTxy5loFVKpAkj
souCojkWXhXK6zuvU6oipNTlbTu1CF1MVQ7GgLTTQPGBhZXsG5cW87WNm9n+duAvm1FnlGvZFJib
bLqeCnbhQZToEWU0G2nLEEE4052fPAjy05xlNNjCtnn6YOhEKB0KDDt2SlE7mUyLDQMT3XeVePJE
/48bYZ6vxm1Rpo0DZb5a7wHAsMO5qoXPswWQITeIkknLsyp/kiOi9UVNvOvl1KcbvEaxDf+C/rNf
O7V/t9cg3sgRSVR4knbHaJbNAhMNgJy+R7NQ3SQflPv/yvlIX3OBFiTszRNc684GF/zEpBumjvmb
I9LCGF/gBKpXUmR0c8FxZlcKfnv2yqmF9SLqDffi6mCiXURttkUn5nUIga/ZCniID+p7awE+wBVu
q+Z/sZOFDIUcSgBHV0ca7tEh/83oguAg47xuMBtKLo6vnTvWs3NJD0BNneZFMtUO8bJ3OB4l2bnP
8i0p7wkXVHhtiy51Vrx1geA+HTad9eqgnP9MTrjbenBADFT6spTydupd7SP7eI2nNAvlSg/YfTyY
Bb2D8myWKISUEmTz2IDuXPpXj46eZc3OZCRusm2EklYgUnGv2vLRwzBtRhdmhmPM6xbQkx1KDNBa
SPKnC5sLhf5hNGzH/OJoV4eV49bnvVvP7qGvuWI6+WyqDGTQPN2efPa2gnK4s64JdZnKwv5oTH/9
Q95Lqw9Aonp0QQNY4ZZ7KUE89Un1Swg0sQ10W7axMTzzTUiAYI38JPMjeqL5ZVCEWBafgGomqXi/
zz3heCm22/GMNvoQ0EoSLcKkTHjT5sWkelSFH4PN5nb20VYQaKWheFz/ycy/RpUW1sX5XtY8Uayv
627tmTuUI7PvOJY4el2T9oZ7ixcd5EpnZR0+UQBV70HRWKf/KoHgLu0uGBXZYwDYjBpvhUZsINnP
GwxBWC7BNh9G387i5KjZ+IPL7xPCZhZhtSAd9txwJkkHI6fIpkPZQBmzKRGd0AJVcIq4UnErN0vJ
RPo3hAdzXQNig/1upY5YKP/IhtkQmG9hi75GlhPBHK0QOU9OaWnDD1nW7/NgfD4d9VEviELcPWJk
oT6g11/2CFNub9yYsr++JNdQv/62RLWLL6lZxJxK7QrYD7zCyygKXHyfaQ7SBLZbBXhX2jlSKhzz
QsLXDlthqz/rD2GYLMZ2vRAwPPyENH9nzmHycaKH9lxKClWrZLPbrDLdUJhqh/zNbKIwa1wy5h2V
hMRK0S7LAjzTDboZjaTbVH4Bxw0iRj6mwlPdBKbfZMZI+S6Y5gUgY1nYsBYvbb0Mam8ti8CeFMF6
4gGnJhnfmWeaLrAOLbW4/5JRWXxpHK209Zvt5Cbqevcv5fdkt3mFqdVoidDfLQUHP3AcjX1pldHP
yvQl/NjtdgsC6dVQbSeZUD7QtBEQlHQ0mcoSTa2YMh/B6+SmF/T53lp6/CgiNrxrFbn29Q209J/l
GVJxCpQvPyRUs0si+3oFqrVBCYDCVzvsLiLPObDOhVm6uOrzYoHkQ/G1Zs9HSxu/E5lLpbRujGJY
Mfn6lpngW2vKRcCiXWr1cBD6jJTGBhD0zVPDxyFNpRCW38DLxz2i12LYkLJm9Oo64dVCvGOPNiul
t234SmTTx8fdFjvYY3PvYLVMCKoowOqfzsr+9KaYkInG3J4znDuEo6qIQizQ8SmzaZY9Lx9dc6U3
CKK61kNxPK/uABOZfotEWW0oNEmdTzQuzOecHzJOZ/DoMTHBdYfSbUN4TIpwoC4pKo4R/rkNbzaH
RAyio823RiHSLea56i88+K0ZOn5zMy6CTswlSzo+OG8VTJOWmlna1nsaJn2/7sXziInOW6m/Xzvv
Ez2pmWpyRtVvKQff25RwPFlnCwpr1XSpdIl4wvks0+rXXhyPDs+mLH70cOEfmLQYtnC0bqOWosSp
7rDe5CB2gXsLubcYEvomBY/DRBbIYtUqFcOOOGnQjk2WdTBQUhYFQRfKTMbHTRZlnlYs/gQewY6N
wMvhIyAvZnldatV6obExXD3VcpEB2dbILTMh3/haj1jAxqGn4gH14bhW6cDRXTYdL6kP/RGuVDHS
FoALRF5EbTPlpDe+Rzwz1AK8vHnfYr4zCmOGnJj/+jwJF8szA90Te0gmREgVnGDYjjBCYan+UL7v
1VvjiltLIGL0n/vd9M30wE2lUN3n+E1DXZHAtIOI/ITaTyvoGb1t+sfuuDSB7kDQ6lsg9pYG7vFY
mtRdyF7cbhclfspghfncoKSPG1lYvhsnvBcnWUfXfPO8UvfUOHYelyZ1xPjV4gB9HjvmfIq9W9LH
gin9zkRbpbd5OXobM/OhzwGjxMXC4XWsRRHbqejVAtu2mVlNkTzBuF0l6C9Da6nUFUI6IGBUP6yM
JCfYv/VBd24twGHUqsaPKm7q2GAauZyZN3/ICMZqdSdwUxJUWdtLQJ9LPa0L8x/XYvXqzOmNjIzK
OaDvPkxKfNMO+hFLc621/WmxRbBU7KEyQDFIFIOiY6Eq4OBlDMD1BavOyKpYwbRxivSQK3wAJrSX
a5jsdDRgBkuRXb7LUvaDOqIrmKXmrVvjod4uxr9bi36WpAzPIF9t7b/oqiEfmoAOjTKSX8AZmWSl
m6DAPRsqZ4IrUwAV8ygQjjWJfDUbWFpDVmiely01UVBfENv9+55oJgu6sgAjX374dL0KU2OEzarv
ZS7lUIX+WUT+QTOcFOGkAZeiKwSGwTQAGAQwkgfzF34MtwrX4iXF8+turyCC18eIYpebcUq5WESN
LDLkgGLJ5DLJlUPfiUpJJoixv17x7MI458AxW2mtdyXI9qm87jwbWUiBJ5dE8c9t0Kmhee8/ADpK
2Aernoufrg9GZFA9vkkSJeRvRBsCIRdVZYevTo3GdDW8gFi5ldeX0N5q98H+azY3+d+WKRLt6dz2
5wBiJTPqrKj1Dnj0/OEBmulawu8V8xeTLgqtqPt7ZRmdTlMXIaFQASAJ0YDzQWoTtdYH6NSQ0F3O
O3EGPX/Wg02CpGXz/fCLICbAcatzwOmqy6d0Ucj6p4UYuwfaHUN59jmNaLOnY781HWn+1d87wQQ7
EhWgDZwjwM78zG+ZLFD21vu3nQIcPAIB+hDFiYJc1PZQwneGiMo6i5e8wbyBqlhn3z7Eh/eUdiw2
0FOZ34TfHY+MK6DxEpmTvnFOAK8hvB5wU688rM6i+cpoc5gEjUc/J+8+QzZ1ysE3mhuNzKHBAWeK
0gYbYf6e/0Uw6Yw9mgb0ACPkbl9d2mBPFI63GqztkIP9gFAKTKXFz6EdU9/9uwAoKwWRVEwyLtmO
2NtfAHUmhxNImmEGWzWftY2qci+/t8glvzI2jSq0Q2TSkHJZpP9z56ZRKTlyNfT03WbpsYsXCw95
0v/dxu4vIO8UUBTbLP39FA14822+CKvPMcqI5pj9elbwAuirs4KmoK2v57QeeYxls4+1c/ygDJ7T
76scw5N7Fu2Wke9eO7ApH3ZzkJGkGCs08UIsE7XKv6eawgRkFhs/A2C5/Q21OtNzsUUMH9tA0blL
dclEnnea7EIiReiNxpuXoZM3MZnG/4vq5CGbyzolCcFXv4LKkqjl7jcl/R24yHaTCw+DFuEhdzTz
PcU7709dRt2tTl5+Nlwrk6QAyf4Gbk7cX/01ZmaEr9LF8ARCGwy4clrKVNsB2t3lJvWBrUjXMUU3
zF9ejWNCtj15h0Tb6XaGCz70P2hIFS/JGBIWLZkrAa+rkm8Fog4t1ynK2hk31YhwjIeZLjYB3bXL
XcvTEXNqwcVa9h2CgYd6sU28Fw6IgWhlAmtI8FGzDC2wJROuxsy1nXHmNIYJ8KoPeNayajIeveWY
TtvV1sdjIcJdonIPHHtWv7k/2sFx4ENHLodDTEKcdYpSufaeLAzLqOriBdqon0dgCerDB/W/zwiX
66BA5uOLMlz0Do2DYr72YKaLLSB3YoZzC/9YfuyLaeSQRKzYkWOy8GRnyFtfSqh673JLvp0efLok
oXekoFp5T642SiL8cXja+tJdUUnhUZn0uauA9XAsRhN/KnMs4QWo5PkheDNM4R3woQgz11ZZ/k/4
J9zBKrwbBjqtt2Q97Tr4ZpWB6DxGotYja4yElQmDDlIMaIeUY3IcRhqeCSWieu6hR/pDEJOPMgYe
JMt5K+SkqOO0yTFCoA5u9jtsUPwbRh+nQD3FPqqrdM9PYwVjbdQXbGuAB3rFP94PgwFxcLyOSCLW
roHRS76sYg6Nu0rehYIidGibcpjlg5Irw74oeAVxEexXhzSsUByj6xEiHNJOJMFabmFCPtGdyXMG
dAAVzCH8VJhQJ2eK9k8lpMFtx4ep/HKFQyIbxg6ml4cAflh2AxjJbIEeuZITMcDPguouzDSF5xRu
hLGx8Lsa7NQXuShH+viizvngTMgBcDvBKZnqMfmJQqXxx/IvXVBlZNYTRuYKvLSHVNZn9HL255kE
Ejbtv+/vZoLxyNcsWEeFNyE1NkMFYg4QwMGN7J7Vhp1vTlmu98J/L8cwKZeRKixKoU47D+4zspfS
lpWc3AHhvo6zijs27iNDzShd/n3mhKkwfJp25sprlIZl5SWw/2h1VKowxDZsizMa/QqxdGtW2x6u
6Ax7LQlYP1Og6Ni56ESzk54wmBxrIQZDAryhEjBPA3s0JPedDTFT2I5CBZfZZnsXbyLtsTOjnLkQ
5VwGOY2fNC46aSupYUogfAAH8wczACYTtcn5Vd+Y/2Zn+bK/OE8wfnPuYOZ8zonVRd0xLnOKiySo
qG02aPgc2KhFn0eJnuqHn5kvgPNRqA/upH2lDqtS6rF85ZzgRriPhc1tZpXCv32/zBmG9K1mSHJF
Cxj3IFnZ+hSJVPELaVQFJbSaQeE4sO8qO7XbGwEmZ54/HksOPCS20UUvhCXpYxG0Y3+h8jzCD2aH
FXjZOYT2hJn3IlUDWOMyuIEzfVBCpAtx7ysk2BTj9/a7BuEFkCF0i872usqC4lc7ACMbBNO3PEm8
3DoxAz7qHoCkxpQsAsbCTaepmdvXSx0dkUQINv1vu84TVP+syWroTJYo47d3yIJVVeRSx/+L5uUu
23E63FO/apx4sGug1ddChbU3EUvvikf1YrHc5+k+zoT7h2tf7G9W+5BJLGRcCX4p0Evr1TzFhLON
VvaP2yE7eLM4LVePXTQdP+p/b4apFwiueB8hP0mfT3b13LJuMBAIwxtDDFaOqfpDQIJxbUV+bdyq
0MW8NfHMrVZKBkZKiUJqb5AXJaBXIw0R1xlK3awMUKxGbqGcd2tPe589vcBDtUS2JqsvMRGoZUJw
Bf5Vns1Szs4I8YXz8HnjHL1bQXArtv7JISdEqWSBYunQbi9TKK/LXDUXmoVj3LAqAGVF67ObEFaA
c1iI6H9iw8Z8Ea28xmcpSPfgzkpq8QIEp/mFJeacHmqC+xC6BVZQZhOS9fIgs5I6WctZDC3ZC4mk
BWgKWzZB2bT1t4+0MkAj+p3Y7RcVgNr/hLAsVVYkMn6GuFLh+EeMtXQakZI1OyMV5+In1PnvgQRV
N3+CIqfAVNR0+kk9pKY1rh0oGxtCSkeRcKbsRp431ocD1PXv6HtSroBqrCBjxGKlyy2uhCEKKxiA
KMWQfL4quhmkxTuC1hOn8MaHonwXBHc/2kc/+yAaaO7VF+aMMLAFJtwjU3HglPJGT88HeEbH6Sc6
xDNMLocioakVVnBV4Iqk0xnrxBAAyaX9eVErOr1Pio+9KaaqdqFV0erhAGkHqwDbrg2pDE0x24pf
YryCqPbxBPmivmNCCIk+qCcpGG+0CabqAoY3sgNAwRVJlCb8qojJvP+wIRAeSwfjrD9dj6E14KEI
yaiEusQuTI91nufgGyASv0wQGfiKn/TCY7CPLDzF32yz5EWc15BkXz6YrD4pj5WcIDTtcadNqSCO
5BwRAha8nBkhcT/2XnnffJCjsFB9JUyPsDptM8fYACr5rrTcJjv1/YXFJrf82j3OFkptkoM+YIFr
fQXB4yuwQ/b4+3t9PslqShcH6ndGmbUFQegUGNigRS9NKK9ddMXaG80uPFz3woghWTVovddYxaHt
NsArO2hFYcn+m4uiI/KSeKMM/aqfIWywAOZAF/iEccRqIcFw2eeV7Kh2O6GFBzpHSUaNqKPOd1aS
QxpSC1BtmGtltyrqPskn4340ZDuWPMl7q660kE/lIAXphzIcdBfREYLTVfO5RWxgRdmoib1sqYz3
8dwH1W//4Pc2yHchKf/60rp7FGqoTslW8jnXrnKWQ2A82CxGgNivH1tiW6XCxYagOF9kmZZbVxWX
M5fQ7g3d+XcNJi1HWnWR1rUa5M129JWr5OIC0httZ/0Xcdg/Y29bEurRTElUxbavEynrHdLSAU40
DTUHMB2+I3kZgpnwAOvlOOyCYbRLEyADlwnplggqRFQ6Uuzcdrz09OVm/VdWlWIKzcDWGkDV+E4c
gNscN7na9b6QEKKrSSvCgRqfoqkcrTK4nvOH/NvxgLK/OP6zzjPzmOEirJml9gL8MuqDVEBoZkG7
ZypU53GmhFnl0KF5MQZ+FO86afzb+PBA6JEPDdRFhUT4O1oRKUYlMmfs07+9wnhdYZx/YBvMW92H
YROJNtddR80jsAUCxNOvPdUUVzTnSoo08h+iaG4MNAUBzZAtty0pUSLzELHqNo07ReF7cII2IbrH
r2SXPt96F2iboTedtFyOHLZgUZhpTYPP1R+l4Cyk6fB1Y56isf7yFgz12rL/JE+5GzJiL9TmjmNz
CXedT0UfGarkG0n3ycmnx4AktcOOEl9Id20pnrVEmJ2BXa3Vu2hPD32rGWseSyTLAsvQb4Pu5kZq
eE4MwfE4gqKuO+02ofL3IavQgOhhj1oVdeI6iNMbrLe74wvHSXmZox1weIa2yvGocIL22ghUHUZ4
pv4FwGOsZIIJpW5jrTYLe3sTdB5MhVFJ8eBNKU6iGSPLsUiqiYpOLCg3hHfzTqJMvUUQPyQcewVu
1MJMruCUhF+uhgW9i9lbIHX/1eTV1TC62MLxl1eI+i9IZosqLbhHtUkd08gFv39/ngvM7u1hfkEU
rVqBkWNQrXGoX7gaq/yxP/+ujLdDXnQgkho9FmS4/lV3QcHx59Tbb8XPgwfiDYIOB1Ykc62pDb9l
a+JpAti4sKlxceuxl27xfD8gsCbydtU0uv3klw9LNGee+ej4boXvDFkErSkB6U1X51nIj6v9pywP
8H+dJAX9gqzriYxj3RBqGprvPbT9oQC4JpLRmPl291IsO+308X5xhRvm+f8edlFruLGfBxheWcvv
rDg6/DB6Dx1PRLP2xP6H07pWi68ELKuhT3rNOvRJZhJUksSWSBP3MdUfEnxKSOM1LVhKpEg/MIiM
GP55HY5Bb7OR6G2UyK+sGXbIobx0Tub0+/P25ZrrUbubC8byVz1sF6D2wIhMTpZ9Ht4vxZu3IzSQ
8GKmHbPLUmsG3GvAi0KO/1KurIcjoTOmXbq/fTSc6ENMtCDXJ7JkfRCAzbz3FXOytBre7JuvAPCF
qN3EaqSTBROHj9VuQa8OMeD+vEFlQ07LvJFmbBHoJj03v1q+ztuGDNEzS7NS+BXOHXlDgIPIzR0Y
Taubxq9h7NQP/9BJpUUuoFGSmIAX5mC8Y5kvF7v49VbJtHqQbUZ20kWdPcKudWH5q5rFUrPYKkGO
lfFOR+Csq2lbjESFYJoYUecp26Mt3XCQ8if5s1lSQVJxBxeREh0rWNGoxckmMjV9VGpRsicfoVWd
fRVdeBsZD4/toMb6FrZI9pKOA6wReFHiYZWdAOLnfY9RSoJ3B/8FQ/uwmPhGlLCXcgzt/ry3/oCV
1fgmm3qAbas0pkXJ9kDuUjANjmHTgf34TstzcnG8gI4jN6TT6biy262H8dNAE4hRQDM2MDJjMPhV
gSXrtvgcsI6+1yUItybg7eaANCVghtT2c5pLhGmrywIbr9h58Y/fjnWNa7aOA1G2Iibb/B0KVvyh
I6JtZKgdlm/06zx7gt9R3nV104OZI2QiAZm+Z3Q5Wp1pddaL7zUvtLEvPoYQLKvaVGO0dWAR6ljx
wo/bw5jfvU5k8aQ8iBQ9j/oP/mtOVSuaOg855DJ8070S3bQGEbyDRzIj285dEv1r4eJVJpXRoe6x
ygKLUrwHVoegtwfDmh2mQ42CszG2RKnbb22AUV3CjnMgajJeaZPze3Urz18k3Okscbg4GFg7CJSM
tejANmKYvKTsFLp7Bg6nTo7OmEYZHgIKka8/nfXLltRBKpSpLxoVHSaDhP6RncxGvD9hf9cWhKUI
WmEFr6ZmmmlM1IJVgMBIFny2/CFBL6GsaLkupvBIoWWxtI9boISgs+mZUuW6ad/Sq5xPDRPU4niE
/j4Pu2SrIKcOEc6a4OzSftruvt/q1o4HdJzMqBWn3Xy2Nx6i8UhG0tyqiJhbbTwLhdr2bAtDWpgQ
iDFYUtqFlNGZNZgNBAx/7gNxGgW2ROWabossngqt1WR6fcwQV2IVYEskutd3R6f2g1oWJ+IRK81T
M7S2vQklJIw429mX7E8JrybGN9XAbXd/v1hOTfpKgKBYxYIh1p2P+LySLTyu3zFk0wIiZ8Ki6gos
TKxmsRdILo3p2rktQgLkMJJ3n/GC4lXd9HyIy7MobMb3ovrRQJ3l1VPLZ4UgwsE7iaY/qkpZPX2L
tMPclfzX3Z72wB/LrymXSvTBY/KPjx/bR4xVdoxq4sMsxBYlz7h1WJv8350LDAm03XVGnPgtcaxh
roETtNf4ePCfKyPPqB+hRYZJAt8tCbcnrhebewOe+GhTMO4Y/PPQDGqfcvjs+11a5TOoxKfErTId
UJfyQ+564yCO4CWq5aCUwx5Yoe7i32SkWmKKH2h2DIJlv93IcvQ8ydEYNALn/d1NcBvSwsAHmuwd
SDzpeOghym7R2ISTa7tKV3rTEZ2fpVfpq6TiviI5MonLegNuOj8ye6TBSItsjFkZhjqnozihd4Kp
eWjPUi05y4j8ax8imqb4hswEzRGcqZyObbVsUuBnLLS+8/WD78CDns3iL9r1qbcH87Df8Lsy2oEc
AfRVTqDpa/pfp7iS4Hi22vLF/77qh58NYCAs5RIJBQWK77PpFsUGJ73OX0S3bXvk4KBj1XB/dANS
ncTypD9apk+RAvzG5a3MXoCErvaWhYV4Hj3j88FdI6TFsanwrhRwCTX1QGWHRnAnh037ctJzsuAA
kubAdNg9Km9r+JzZuJQyVcKitKOH8i6KeTkDZRxJ7/oNyVbYY0NEHFzoOpj9USbOomOYPKJh/MQn
XIP6r5TSQxIpXlOqf+ZygXfJyagamjwxSvca8feDeZfY0OmBZE4qd4BaoGBdkCs5UX2VO3pKpJnK
p5ynqcjPaqR+1b+qWkuJoDNTM5pSBjRFUfzFSsF7dNEnsL4hPse3QtfgqoDX1BbrK1XLFdOok9hT
z7IWoxQAYT6im9rCVS/mc9s2ABhJUHY3xR1Ls7Vkk3uULgDXnlmpychLA47dk/GYsHeis4fhVRIk
i6TCH3NjUyicP/hkYBkaryhTGMpJ24UjaHNVQjswC+sF9HiHfDzFkbIN5focJ+i5sOnIgJocbb9H
dclctrxv8MWaP1QwwjEVj0TaQ7IMPhbh5ZJdyVsTX97cFx8iL8UF/El9JduIom+IzxsS5LrnZwl2
cdzWFmPT6iaBOfLDFK2MFoPoNvmmmQQ9ociG4E6J2s07lt/L5/j8dPkd/Do/HRSPS1wFBCilHurm
5hxTTyOMAZ2Z0OvMPrIFNs/lMrWTDbzEO3T1uEgWsunKb6D+o6756fAdCASAzsH99WXZngEu0DlZ
URAFgJ+hCRDxpPuhzBH+p7qWek+K34cKqRcennvY1Yj7KSeFkDgdEwLbLx12++rrn+x2+3HCDdNU
4/z7dfnSr1eX6SOaGoz6/RrrrMLjVQnd+8RzY19easjnxyWe+AecJF1XF4187nnU5cE1R8+RkYo6
Z3gRLYMDG4rVf9p+ANj8tsjKLOXI3H/wd1xkXCBUvCIidyIyEbjUKHeD6Zy9Q29LToZArmmlIRip
w26vCdXnn9cOLvvd1iSPvyvyVk03KvazzNHh0n0eSeISK+QqUuOxuyerX4FJL2JT/wPNjoS9yweB
xpHyBdKXOMVBYGcD5EfnzrmOOGwtblfNngSvEBL31OU3CoamFcQalFNZ++EWYwXjTslIVoPTB6CG
edup32jnBnOJv60rfAmVtr0x38tk4Zmj4Owhcms+aY+x05CRn3UwFHbCHl5qV2v1BT/WbB5W2zVr
fgZssJKspX1ZCtL/xZxUm5iveSUY06Fk/0+N31WXuUl9EGij8v8sHnAH7bVCgpeu9444CbtJb4kj
H7GwqJ3S+ZaXZ3x1k1UheVSoMi+imMWw1fYTWna2PvwvPz2HNwgPQyUzyovM77DbZ369dwvo118c
8dW6B1lPiluABDqKXagPKYCwJaZlRCGCgYoXSQDB8GRwoyDcgc0iEYiEdsu2tUxJp+GrEnZtBt2O
owTq9P+7Yx2/tEoYjmuIPFm1wkVbHX34+l3LfROHG6OTueSlS91lFAOQcxtzKbuoqhox5HX8+a7I
E59nQDQJCONTFmutAMCYEc5yHRaeuns8Xs5OvJvsedfk1PnwrkOlSSR7c6BzWgCxXZJv1aRw5dJH
sz1umMiljnZthPpTnSsrgEs9KHOxAEAs5RlzMV67mjXyaEr0Hzl5RBnuoNXDpQIcvsxonzog2Sko
7I3JuRS9lGW0kC686UZgtK6Jk7fAFdzE1I8+e80weVCyCmP5MHs4NJE4boXh0pW+/kLh2M8Zy0EV
9avDgw6tAZFSAQ5+yUmsjcfMY8dL/eWojHGuwYTO0T6Yjb+kyfkOLPaYZMXq/Ehtqzy+0ZEhfQMB
6aWCIzp4tByNhgzXOozDKDnG5H0h4KCINqt0LjpOkEA7L8hQdb3+pcOxyNBM1lrICFWFgloV7+vS
qFCdXAybIC0c2gVDnwxv2yRb9zEss/GyC1CyH4oBqbSWGlCKOzIeAjxu4yMJuiz4LA1Cmbw70eYF
a/Y11JAiqjl/slTWpWwhSWec/qZszuN6fNOZuxLGBu+R3uBfyQ0DWPazZVjQKQ0KwF5DZQfJ6ZiH
j52TVsL0Hst6fZvXnzQwqY2WrTnow0G0wCFKNlgq6FrhyeMs/DTch4YCg5QoKSR9cgekiZ37SF3A
1ULxTR3qYxTX7JnjHAV1QdRKMTylivgvMprMfIpMbGk9utJm2PYi19sfpj6fO1IoBkmzyi012xHd
3U+vsIFlLr1ciMuMiVPz+cVFpe1JYYMMCKfDqknQ+3S638jTESzYfIwKwUlVXVs326LSNXdfKZYQ
2bhKA2Y0Fsa2YKt9h/kCIF6TbXJcSIt903hxiBC+++dezGKbs+xj7xuSTwoJYf3WoiFRmF5p4zJA
e4My4X1VOsZmA4E7QGPW9P2/ZYP/2FCMs/78f7lydvRtpZTDaRjMEKJ9cMmOgYnxLYkNLFAhE+bs
hcJaiIrLkv58wJOdDJprAXuOeI1S3jDPo1Y20jrdqE4gZORzKjGEOgQ0bi2+MLgqYSKfhwZOpsCe
M09rhSltNJ/rV0SES0wFx+dd84VLCUK5bCYtO/izL3+GNpSPmkGkv1KkVRg6CRFmDvA9FrcenM3X
E6NDipxt4nxr6xj7RlNSHbJIpoMTuKoB6YyEugfIjxFs82PLB6RHGRRRflewDoRmsFAey9jtV5vw
dcm84xyou4b1e3nw9/gs0zUoVnbRKJRbhtx8jW4I4HbZq4AO0rCzy0QzQ1mvA9Odh3aWWF4ofbOf
7AUI+xqkGfykU2iYKyWjcnPHHJfYk3CEvP8+V7y6+d4mnw87aKOPFpUsaQFVXFPvH5dM6kvRTLp7
6Vc8Py631liD7WhI48qVZu8U1hc8H7ssg2sES3ABxn4yT0o6GW+DYIZRvl2ez8VZUkWq13c/YCSR
g6te+wnpUVSvfm5+SAtMe62SEiiO75e1yHmG7dsqo+P3eHmKoRZwjc668LjrzNFLk2rntCl7tt3E
PawPXfYNVV0FRO/N7eaMOVZ9+D3xxsC8ei9wAU8Dj7RfOGkycOMwaaFkJwBIgiPoWt48FZp3hDgY
gtgN4djfJkhBxk2IRcFkC20SUSPzSSiVKFB1K/WgaUhy5AgXhQs/1yeer6sMqO3A/BMAZQQDwIpr
WokQ5MREQdoltPuekH6QNcale19fbzpXV+zCJEqb9IIfrJ/so2Lr8uLa2D0b6kS1Y/AzYRlbdinX
uqV0h9TimH7k5I5Ued/tPoe83QTjLu0LO+KNYLA1HlJDm5nttGCU9qNWkYHykaJpWTUgsjQhal6w
RfJXbD8qbuLqu4xR0RjXzP42DzMA9Zd0VJFUYYsYBIiLqYJw4yL27HdjkS90BzBiXfou2C+Jt7Rm
FMdqH3bEKfdLxg8T7scXdzmR+nmqAM8VnSEZZluEpgKScxkQIrYg3Q3vFegca0QdQv4XSfBeZdyI
RUjVTe9dby0lqK5dmsszN7vHC+/lpBzdL/nzcfvi3OyzhWXeoF2YtaeisvyI0weuZTGYz2Yf6sm2
dkF9LxTK0XJX1cdmuZ0Ujv5pBfUYi4xgxayIJoBroVdYm1wXiS/s/KAXoKEQm3Q/yFMLP0soYCY8
z1dOlBzLW6kHZpR2+++ljNILuuJJhXzZuHRLY9xEBcaTrwZd+QwlxOTCwzr+xPQPqiY1RRwpTrxa
ycOeepBJQO3xCL1WgH0sVK9NeYzSOHW7Vy1ukdXoYCCXcRig9EIyUT4WcEIPKm9zgqgfOMau3OaX
6Ln19eXNVheZk7S9JAZj8QyTlH95cWmUSb4Bypada9i6Tj86nqr+LlRtfAFAYM/GkZdZ/oji7bQG
RM917sTxJbY3yhwe6DVonZTiN1d0uyvEQqzSRPfdLY6R1JM8/ojlh4THb3hY4cFbB1Gkp+IBT/L2
sACMhWQJNZLHWHxFvTJWX4hOpxg9T4BHpKK3ai+RNQYNIlCgm+g8RNtNPimTuQW6JehaoCLv81PN
Aukm9pPXeF62N/N8sJ8mxd0sqwNza+dGnYJ1Ii+jXyaVSK6dcbj2sagllclzbBQsSrJeOq0IGsoT
yWyQLaZ8+2Zg8gYGw7p13TurTfbHUr//UJqyeVSDLNSO1BJCKuY0VaXZQqfSYe05jm5j80ubAsDQ
Ytm0/G2i/uA+quvhhb87cRoLFOirNjU24RMVVPhGTugrBpFy2y9RdxwR1B1yH57VGfLXmvmWJZ96
CG4qTEUfn+svbV5MZgmOq+8URTRJ4+7yXWR9hKpIcxDZAR9zpwDIaDqIpL7TNIkvdYj9CMeSuHrB
Qm3SIlmV3PA4CWUtkE7rRLL7AEGIXtRsbM9D3ilFry9FpMevZuEtA59iGELB/eznuTDqHtchzTvj
I60I/57RcnC7p0ODzO7aF8lofNogkJJkKEWts9hDDKSotv+6fZ5Z6M0ADHwJz0XVrBhGyJpu9wLT
pCo8BAJ3+0qWN5YC11fTuuV3T48rlCLxEg621pYkYBKJzfH10GMlHoBIDfU1y4q5G5PVhJOY+hXi
3jEWrgPnuHAw/VVnMnYDzr1Tb4eE9iBowTrrgK5pze4vH1nD7HYcBMpGUKMr4iz7ZZA3Ecv9azN9
bXCYXz2yZnQp/0HwYdlFuJPaqT5HclU6VtWnxV3qgIJwG/WKbsdcXPhjYKUKPwhSqVEXRnX4Om+b
0x3T7yivQZFi2lOBVlMQprlwuRHIjV80sfmeso3RvmF9fhpJqf0uLMLZmqNVHb5C2tN7QrGEKQjN
7LHTiNWouslciuxeYSbhfP+q9/QhW9Yr9INhsR5/zVLI3lfFu/SU1GBjFzsjQEq3WaqyGKQoHhzx
sdtqGF3fRP3d2pOmh5f/qDuAWUTnLhXDb288JyoG0MrFTxIIAv7eAmLhdrP+yzR7NS3HUB1cshgc
49lN/kRJB68A8YWt1pshayO2Vj8TAiwBdnNqxSbMcZfoKFzgTNMpDQKz2hSFro79CJZVCHhB7LF7
UB7ealIgN7IMQvTNlW9IGiqSjqISar6C2EzWdjg3B6Q6njwzxtI+R0wyd7VvLCqE/jMdfjyiy/NG
pL6v2gamN7sa5cx0FaMvF4DMqrOLUMjFLwh+RXtb9jvNXePmhweNjZKy+gm+8lnzMHU6TLefSKf3
4wDfTiTmHvhMShhht8ykJN5qL0Cr8mYLJKZSRsksafW0y0JIzS3zEx2CVOWcoRifehwishM48cVQ
7FqUnouia+i3K8ZxajMnH9lNL4nDnBplp0HMk9pDYEcGwc15PJzZHidbX5byuSUqbOn6kcOY9Jpi
cpaMJLiJ/zzyejH0CwE8ZYnAuZ0eskoffuvlWjVyy+ZKocaTjcj0uWhnw9Jqdsnkmh97NjgM0UB2
1Fge4NPNfV+CdvHFVOyaWnU1ns5jkQk79oJpBqzYm+FpniALCvp4EZDToKDF1r732eyopekS9IaQ
T9FosKaMOXuHpIc/IKNNwlbtLkAjqPBF62zRXcjpVH8XeLwmn3rIb0W8+VKRyKDnRNUrCqh+O+6Z
B5DxnVpXkcCllN8R12uwfkJ0IKZM4YC16MeIoJC1c7vq4NvpqFUOHXPGRRxIWKIpsiNGcE3vyN3x
W5lZCZNj9WYFoqrRliXAvLPFMz4teOiWDy3HNJPt1q5hrE9Z3ecEWxgmwaRuFVtlJb+WSgYXXjNZ
5KP6QQtdj2z6JUBUzsgkAQiSDkkiifhlrRY9i2MP4hvuhHkL40hYsaFVCsKqH8Us4h6zDtULEkxy
5S6xKCA/I+ZkkLlLaxRAtL31x1tIqYoKaZX4CKixSl40YipKNy3roB/Mj5wKUSX0/g8xtr2cDaZz
TeIjc5wC4yy0pa9W99pRfFCKQQedWtRTxH+7lpSd8YxC9Axtwl7mHCSmjpbI2HjlzDcOBKRsOcLK
EgKI328CjF04uJ5iqyO8PVP1WBqzsUgAybdtVhiJUGXmjOowJlZTn9vQ5KAMKR5nGL8rNsTZ77L6
rj/duwoVR3xAtpshr1/o7eQCGPBAS+kRD/jJM2+W96XgDsKNbqiXlxaiNzlOcGB4/ng17of6ZZ+O
ey4eaiQmJlqECVIy33NH38Q4a1mbd7R+dnivKEm6IsxGuG98jtCNVuIOHvWMVrmtpCNtmtLfZQx9
Izyi+tXXpiPvlIyvb+fmZ/5wA23KJONBopAJaZVIn8sGh9Xm3SmpDnATB3850ZfamJrGHScMxdHc
J8OgAZF1y5TONq0wxL/ReSxXXoxay/lIJSB6jOB4yWM9hZHfNFPutk2sYprXATtrPmLIeV+PdoGF
Ee1jDn0GLNnisLM9ONECrHxnRkn33n8Vi5mSbLF7qorLpEnkxP6gUeo5CDeDRU9T7of9peWmvH1f
shcJnA4Pt5kPj1T10V7YY6r9ZbhyVAi7E7dbfEy5NCJK/k1a6wOaKaQnzZurmsAnWIN7rVTl/vAS
mGyryE++/xlHu5deEjQ8llDSyQhYa72n63NtbHzMHk4vgFnrFMl0S5vV7ZU8n4TF38SkhTuYXbaE
SIXU3YtDwjIHpimo7ZxoqiJyrCtOnIY+l9QJrqQFtrsIGP2M8xeZjkzbG/QYo2KX9c4bQOINBzIZ
RBHoff4SF6znpeRkvnxUYoGV+fATmFWBAJytI8DEeAIWoDKrdwRXr2s7LFezq+tZ+9xkzqqisBEL
7LpmDgNpqcw7C0AqB37hjn5R1HG7LGpQhyR2PPSe+MAgyKP8VvEc1zxNaHXBvgKRXHpmIITckmeH
JxMYY2oiV+X5qTu6v+LS0bbWt8qA4ZqT9eG5W/IPvBmV+XMk7gLqfvUMXLmigZaMihjBHEDL6bsi
dFE/ddc0fnExiU6sfQeQ5hmT5WFGtJwxo48Q0Ja74dpGp0/Cfff8Zeviu//dQ81Rm17x7aU4Pxnr
x3fv5dr1tN7xocMBJNQFkP2/BR9T6y2/zPrRpWOTj+AglctfMn1no2JarWAF3IqKHU+tr0jE198e
aFaqilENuAvzh2JRdh5vwoy43G/uOrx3MdYc06VbkAIbjVkgOImByAR4hwzTSwJMFwgorO/22L30
kdDLMseqf9l/Q6fndW9G1jwlFxS8POu8MDC8kT54cp2u8RPBwPGcsbAyMmu6vD0cc569Jtq4E0NW
M0ZlZruhrDsQSPer1M0a4rjbB/nyNjZnMbfuB2K8Ltu573uaYn0D5/Cn0m9qRFgAt7XCC7enRrmq
J4njrsb8JnBuHdngs1rxbf1xYWSJKs5z5ddWclTLgqTn/eBnlyoVafGiYL1712rdnSCxQsw0YvRI
lLAnC2PTmJdL4V/0txhtNnUm9mG+a1pPFKSaqaxa420jpTd4yhW0rPNyS4JRni3MU3wl3+DJBN7C
oyeXiochqqIS0BdfwYX/ue8dPnQWabw+rnp9xq6boWvsXCsk+BYK7EKUeME6GBRg2fif5srHighA
7m6rP44F5/+w8VEMHqDjeHprpB+OyqJVej9QmW6mKvZJMHndSIEJfTjVgFurK42aAGS7atajZ4zc
TxGvBDMUngEA2PANo0QwQxJVM4RTFQoFcTzqfTSZI2R/9bAJ+43WvWLBWydDOQyfjMTEfXZ4DkqV
+a8deLAZ/IMTsXXYQs44/2kBO2CBp+mdt9zXptthVDXzhG/99Ejv2XRbw/kw03STQGrvJ9XCaJ56
pW1j1vwV5j0vsHoK4daXMk+1k0lsqMFV0wTRKkpgkO0bQSj+/srprr1jKFLB6z/F1xM9dBjIfp/K
Vpu78wvfZP6Si2WBL2fdf0fsn/mh+Q+0SBF3shvUDP82hA6KY00YkAGu4IT9PBsAM/OJHBbaNSUi
5h9Z/gBJYRFKY71inxaep5oSo4hTw5NIqX+tWK567W74TskkakEfnCzB25Yu5s0CGv0bkSAl5Nss
LXSfEnN1sk+KEpIYpqA/T4bQrOiF/Yc9EGatPpGNPhDI+jmY7Ckww/QZ0KoiA7N5UmJTm3u3A0yE
F7N29Ihyz6uSaHhr7/VxmnE1hsaN4Gobm3Xh4LEf2+P1n8QqswsaYSi6jbDLpicJDyqTGrza5Zpd
fTvWM2HjkjNgUNshY4Vut5xBd48W0gTi3hTKURPWAVmkosAq2X5car0n7Dj8m8y83KRsHSM8uXlU
K+6Ash9MObSP1qC/LrfEw1QaRf5jA2btmfeioPdxpyy9c6dYrN01are16l9ygwKsbVDdfB9pYXrR
sh0f/CZ3A1plxN1qQ5Wo3re8Tj7gjfZzajbYwimR6Ty2oUAgN5GJmizeeURWd/qj45NEmInd95OK
VfaKZ+gYCNLhbQmRyahTuSb2c1THBULmpq68S7hn8AYGDf5MaltQO4DwiTuYySxmckV0W+8CYVXH
jtAO9DcrOu8k84WxfrDTPakn2dDs5kK/7j3lC957YZP2d//N2YxLwYLuegrEOoKyPXVHcxYSY5c0
t23ASeDaZgILY2bLD/g2t2I9QNkbln2HN/KMcQs/ui10PttK2bvFFL6wXQOALAtOBnE9rrsMftTR
fezVmqt3ocoXSlgzg4N3i+qLAmYylqASAj3GiwMx8f5XtFe1kcwOJGcFGGIK6q5GyJ44IqB+XFCE
MTqdUY9Mw9boteO/6PU77H+0+obfN1fwyLbpt8Usq3LFhsIz7W0YhFxeeG9Ej1N1o1teqEVGjw3O
y2C6GsyrfniwM1EJ3jh6ZOKwwiiFuYN+aPtEZbylQPUGqNcpH7fc8g4rqSoOAZuWSCEoB5s9+8AR
n0meWxS8aFJ23kDZeFrrQpw4ajZxBjUYY8hzMnWI4OVkUlN7Uj4NOjOGL+rclWVUeASjUcrHvYKK
uM5mDc7ryiP5QD77hCH3iSiHL4vg4J3+k0OBYEpiJAIZJ0szewILotIODHonHckUOaN4uUv1gV3R
zlGfX4owJs5NI1M0hLu4xJhkPlmtB6deYm8ieqxYbzrmKP2tDOCuXwTGxLkyEyPzIMXDo/8RTYqh
O6M0IrgJhGZElVFttutxhtE3tl6q08BnzsX8eHrDXm3AkVsf8u1MDHQ3TmNYjyX1wI2KWsMlPTbO
aLMgmdWuNlqUNdM19CCyyd2o4fdi8vmavBr3Zv7a5o1a25WA/cEM2BUjKOQ7tqP6/dEuvRnCoMbP
DhagGCY9rjYqPJktR2R5iEGnGoA2poMWBdYSTJQ0dn/XK1YyzCv7WcB7akj1b8yjRoAGJWJlSXOm
c+i2F1IJdWNeiNzLAwjJ+3RxNgznCGeF2G6Gl8ZWKDfMd3EaWUG+riTtq3VkD6JEKZEh9IPkjIGC
CxZdPjLpqMCRn3V00ZmymMf9v2ClIxm3w2UAntWvM+ewAnaQ7ObfZZn1Ra4+DUQasoHrv0DXjkXx
VloqHCAEEBntecSC+cbwGg9c8LSQMAexrNLMrwubn4u9du1RDPdyoEhCWGPURvRtuaP8lPNBtifB
BWGPy4id+8+Kf5SQ4dx/D+zvACG0RBb141wqWguTCWSXu1V9GQplbXrS28EQk7lAE9WRM95JZw8n
X9yAYOU4+iND3MxeIqnbkLQXXep3mTaI8eyDQJBE+DtfRmTXW8a8e7MsBOLkjJJnTCzKffh3FxCh
UunAsT0dNGJWVyBxVyQGxbfNUOYawSIYccnVN+O6qywa4GZnvyoaYt+2nGzIv0nfUZYq95kFDvvw
sljzYUt4W2utPiOulm7aRELlHdTCYnv8FUeEBWbV5zqCJtJoJ71kMQkkou1hZuBDJnyIxwu5YJ67
sfWO8/oeXNKdDTAUQ2K2UmmWGXPdBz2NwnPPqrJT5GxaoK2in9HVyLRwHZP8Hj0nR+Ije2XGSZbq
qYrlYhct2aDBdSD6tWZoPEq1uEPlsH0C4VmMnfwsHiALhPzwg6XBTwO54LmBWHOo0LGIUtohErGj
mBmNr3aHGFaCT6kSeEvuVhB/2uEjB71I/dgoezJkJNKaYcxGn6oaNoYR8/kStIBtjGWZNRdoSBrg
Bq1nzpjBfrpbmeIxOR6eysXWPAC8XS5TrBwshOdpDaIKJGfzcSjizZU5scCjf9uiHskVKlWKcyqn
A3wZsw+6sjMflgCDZwgHDXmUdmtgoJ4BnQF3RdkiN5TRp1uLwBA6uxm7jG5NcrDcyMy/QQG6QVtY
BTYKNnuH+dL9k1gLu6cqepEaEGh2GIUJsOA0/7a1Okmx0+wJl64w9X1GpvXbJw35fSqzP9yJYD8f
q8Jnyw5ojDUW1eNayXcRdtBRefzMAF4kv3NAOduI+9Y09/aaFGd7D7WoBNwpF1zo6WNHmpyedb23
qYoyohtfiasB50iohGdk9oncDjRDb/PsFpmCrI3kBaWOPcieVKs2Uuqy8lyBH6pLpgO5M2+p7enz
YzyjV7ZmzrFseKRvlAGJ0OoqPRSXBzBVijjP+7rU573Agf7cfA76cIRpNEdbDjqMDRc/OTG6VJDb
d2SP8gRI96oZ40CERJtLbnCKdqyX17bmeK3QiNKsRAKxPZKcuFHegKTsZJF5h8FA3ybJWc0lEdwx
vHVarJC5iR96TV95IsOO0E2kf0fW5usLnnDXGdtfoUfjlp0Pccqdvh0HC0qpxOf1JSMVZTjocbDV
IgKZrAKcKG2mBVCMONNdvKRDvnsWNbTxMnEKuEJZ0C41eLQ8yZITUqkSB64zIvHGCYualB3pWdo0
uvOxD5nuDO0XWnERvigptqT+WwkDj6fe88fvvItb+/X4ELH5x1HLU+rkMCHeC6oxDF7uUxV9jzaD
o1n7yKxUBocr/q+bFHKxU/XirwBPX9A4Ecz/NOQyxOH9WA0J76etE1GNRwBYTpGgOcUkFTq7GkpC
Wa2eG45rP9gjxJUSeIQtQnWsjuk9nba/v9tphJDRaaZuCA+m+hzqGgNfe7leHf9AuXz0NklXI2Tw
/SsMufaExY7UJKd72WcBZuPAdotsurx/278WF9QQ/TxaS8+0qyUsHZUn7WwIHUKPNRXCadW5aSPt
9yi+UiQujjYoTT/N5Y24KAtKOWoobNQyG8A7Qq++gRHzkKZYN3ECV8mPjepyEZ8wynZ4CJsI6Wi1
1UtKBRrw9Hoki2qY3Ra5cUGon6QUcASIJZpnMgwFxKqI1KcJyZ7nXwNUezRUaIj1rywvzvDZJpRe
xHIgxNWqT4RfctFqxCnudlZ7XpolXdBj8P7ojcVbgv8HN3DGcLRf1beP3pXxACiqNGCT5ew3gtN4
07qMIIoQk+1bSaPqd9ozHIYjGs31zqSWMQWbtRTmC12xs4LowYCjJ8lxPzg3vmg/U/kBX0Yt0DBY
bmVx/I1T1OHejzD/6//S3XfCYjl/nFn5QIN32iSZ38qbZyO3LMhVXabYvs0Oq1JRIkYR9unOPN/j
svv02JRpOOXad7/VoBXEUX2pwqaJPlsKsC703ykNcOLY4A0cE1hS9+/Tpul2Z4kRICAJGlrar3rO
4wlss1ZEIWl/lR/M7cIlX+69x7q3NXf32fL1uNHo6NYeF8lBrR+jAedK3d/hskuGCntJnG7L/HTA
IthM2BT7kSioKpm79lxVKVNVhQW/y8VoynglRED5FoGPtt5vnjn7w+3obplIrANISvvcpWz1vfPZ
vQBrtjTYIyzMUjEBLY5XR5UYILKtq8CuzcAt0nnBSLKr/CeJZIzfiaAgXaPT+hFhOshXei4rr/uw
YtH0dqxZAAKjI/+WvMJC2Sk6J5X+jAyiOfo6oOSQZktU4usVGIPwMACnvIzcPCoFaYPdKiYEGUbB
2Dt79ZKpnMNX6eck2IadeStwOz53pxlGSZuj2dktlwzOwyvJJOgOSvmnmG49WH32JFCwuimkYWhO
Ew1lvkNFAr0qQ8HIyD+gyILNfrFc20nPG/w0rs+UPb15rDjNIfR71+KC8+qAi33jqLkt6KPzecwF
fDzvFGRO2B/AjsZUnYO7NRlwf8Z5QSU6kiLhabM6UkPvODSsSJOzw1o8QJFfcLvsg8a+c0391lWW
i4M9LC/XQ/56/jQZWvnGtFOaH7ppdalbf43+4MW+bj/vRIxgw+sMK31AkBDz77OWBPhu7oZT06YK
9Q8R27fzTod1ONninhBpeKquAZas4wY9XbZT/JRcL7JnqhpVa6MIOX9GeatgmJ1DfLvGWRvnCLZP
XSAfriArsyOtmxcGOkAulLLPxBy5LyOQ6dNXeGOtBxiRmGFMzVt2ueWc58g1KyUi2UsjzoQqDk0j
loL3/6bFsebhPFO1vDQDBY8V9VdnOo6fvSkmDzVEN8dyZx2FKh2mtY4RPO4XCIGboJLnJbeTFU6i
W6bYMo2h7Vu+UeaXkpXgk5/gAajXjHUqR7zAwQ6Nw8crwC8N1QlvKfn9ZcEuM7ENse3dfxAKXVui
4UuNM+cGyWy5AD5qSPKOlotm1+BC3pT7jujsfRIQCrO9xLsjYAKpZo7XmJgUXLSHDPfJNMGgVH6l
28T3O2TbYZDUx8YHGInQvV0VkZKnhz/Aq6FgdJOx8+4jAgx/SoBRXyka4SrJYQxsARqRxAD0kNPt
bZ603LjJVQvSCnFyt1GmlDkv7Oejxjb4T9YTP76izSCHMii5ecjrIKCQfoLlA3D9YrnLl/PJF8dD
JkuY6WZooHS7A3t6KfnYPVPwUysciUQ5mjOfiO9nuRzy78BaFkazc+Heur5QTo/YchiPZX81v6ii
DmbRjt/47/oJOC0AUA5hCHufnSBRBXAXF7+vmLrDHbL77l3ik44N6gXVV5xcPyMS2ItzevvpYtRA
Yqq9hQB3UxVFSUmETj/k6yu64lcySomX0wtuzkACxmmRBzzSro2feew2ylAeBsBR9OcsqD6EKJay
yrAjHnohWdJsG+69Gw+CH3g+uEg3r36RxWeSnnF+WB5Y20z/+3FRJAqgGKbLPM4LFOEq3OmMDCwZ
TcXEuqiqLpqKF7ObQ1EymkvdY0llz/Hdt7YoqtxAA+swqCZBVi9/V62QSyOoNh6C3Iw1Reg6DY0n
4Atq6lE7zCIW1pRTDflbclmigc3SVGWYBg2RKSrN2tu/SYgJACt5Ks9XGHC3RDp/0ZSoHgbEVHAA
FW1pqb0QQ75aNICRZo4g0QGDLnQaVHzV+9I57th7xiZL5EkhhiXYwPcaisfLJWNt4Zdxk/cmR+ak
ElfNxs23XC6c1yX6caxJ+gU/r1DRxjuoXx+DRU/vX2onjgVOpiCANFaz5b76Ul72cQIAWZJjvK6X
1X9owLcbhc5npINirIResi58elkT+muFmC+izcdhcNliDE57YbeUSRvfjl954xZajHQIAyP97TIt
pOSjRpjRM2xyCPFgOA1SBPVXP1HhltDjW3JQD2OL8p4fRUdUhNUrQ3saEFv56nCa+h1/02YRPRbM
X1QyMBIKYe2tkBlr1y+0BXz+NA2YKpl2cAasO4MIPsldA6TBfIH21JGpB8HG/QUpyahvfvXCl/Rh
pKt/Js95HO6YVMxUelNHoGYRixo4D9/FzedVOeuHff3s0eSv/6xa7KzORkxIQMPef1AoX1S52EpJ
mosVX6KtGNHxnX6180DIdL+kwlcJgnpucjr9sJhe4RfFJGqPfUc3cMD8kvA8HWUXCxxbd4QHePNq
XxkIYDi+VF3W29Dd14LUrtbxA6lh7VsQ49HQhScnE+GiEg6P74I+DCQ8IYDbxO8fE3/P8qIz2FEd
dTGVvV4NE1D7SQZo6RS1VVJp7fCiPrnSjcSofZ0fZOgAs1G13Ia26tdgYASK2krxqPX7hr2GljfB
HIlUZsVe42xUgt0Vvw8yBIai3lnFEkCFbaEcjM+t+FbnARy8cbbhNEhnyn6Lwsy4pUoh9dZIh24k
KAlZD3NgLHLGZujRtBYNhlyGKbiAV9R+ZsxFd8tMT4+/Mf8zAJuronCh43sjAXoneFmUe9bdgceU
ViNO486erhPl/Db0UfTNEs1ZLSO7lu5vwYXJ+IfHlo4uzFC5oyopu5P0nsv3rAsjVOq/AzPj8/S0
/HHUvJ0W5rKA2AH1o3fFm7vPmWB2BsZ7lCzv94gUXaUH4C3wbWvro7rq+AaFogEgMoE3pERvXOHN
x9mANKk2VT3ERUMjIG8M6cP6QCioVmv1x5QjnaBFdfRPCbvOX3azFO5qFuPuc+xBsftjDUGY+sda
xvE0jeX1uBG22ND3hM/6KZV4XX5vYY03Boy7OAJzC4p6iSVcym8j26lgSELemAVrfVKf4FAWNYb1
XW8xaYEV1Yh0Zi5IKa4mvvYiOdBhiZ8t2FxZBNi9yS1MboJ/sXHVW7ehu8tmFSCqPB4lDIPStGGo
oGNGdSWXherIgRxHYPEyIZi9nDoGGJeckr7U9SJ/L/uKbgeqQmnobGHjhdUrCPD1x17akJXOv4XB
wfriesw6ByNxVimyNGIO1dRuWCxLBRu6N/QuY9PuuzSRay+2JEHaXkFy15/TNycl+OtJOWndCMu2
TqWHzLEAjSwmkqxM8AVi9Jf8r7VYKKWkfcMxRl919sbmQ0jRwZGHDqTYWulj7rfvRt5IlDu+0Nor
t5r+EzHEuBnb2tx/hPj23zsFZyyMaEh7z7saYgULIY/qWis2K6GqfL0g24vEAd79AWD4eC1wC4wN
r+KQXPOKqYAjTGfW8cde784oRlOLlk5ycD4HvwMnmlaElrtqh/MeBYyHaT8N1HL4QT1sv3YNg7Jm
dwMGomDfuYCQSYBCAMCsUR7DaRO9z4JPgP8PnH9EVx+aJkZF+ldEWYBZgku2cWFjX7wmdmPwi6EN
QnybL7uDzTh4DtP/5pre4U/Iujy/sEfNcdvOAZH9HZz3vRI+NV0TkD5TfKV5GUSChqlJnXeaFPew
6WaMwlY1OB6BRY0zQA4DPv6yC97sCYvV0A3ulD8gEvm07/xdAl579Aia8xnOlCPdPY6yJaKDdZxE
7IT10f9WCSfZkUxVk5dHrDDYnyl4kESh3YoW3I72npVVKG8E84PGbSJBweQDN+6kAqTMbBCmpE0s
zyzfg+thHPQeOy1J5KIpgwNG3MCTaT6CrkNzu1XE+IrGMWQbgf+z+b9i9pMvsWPn/o1LcaZUUIKE
9h6Gb4MUXfx1GVlh3DX5X89d4O24FjZaW7ggI0fdPPMvT1ZuRLV/znz94+MbK5L80pLCd+kOFEAS
dPXQ/9VwWQVhX5M6Ngyr0sNZH6aI1HEHNPr8LC7KyHscZ2kiQfl25d/tzeCkjI78gUWQPntlEAPg
k2eHeLK1dXavfVHXpDoSr+j5IoWw/2mK5Xqp/ayZtRYRcg4mMY0XeKClMPraqRW4ML96E3XmkC6p
g7MFgaclK2VH6Z/5/2bHIusx+wuAarXLRuR5M3POIQ69/P3XuI4W1L2c9rtEB/mXjFtRoWu/T9N9
jzwVSj/fhuS76K8Ys/VCERD6vhjaf8mgqeuHW/2yi7l1Ch4zkqqt+6ptNqFgJ197ZmEpt5k2BvSN
zl/V8nc7182Z3Sd6g8IrB2Ilq5662t2AI30HDTU6QHz5jLjhCPzBhKlgvh8WdHhBWtrzoNpHtHsP
KbeBRh8YbuShKC1lXp4BidYEKZSOj6tmfrGr6m1p8rvcQ/aWb9Kmf7k7jxY7Cmw3dJ5+ocJ04yUD
yu09oTZwosyWCD3be/GvGzuivhQb5VLw7FTo/F5tYLpF0+86dy9a8qIiST5Jy1J+YHfgePDGjvXQ
cfSBhQUXjU0vrHdt8NA3Wy9dbIuQkSsX0IurEpbOEKtjrKpZLzpdhjlUOVrcwDnpONw+VMddSV4N
0mdhxczGSBtgX4F7DfFMddUTXvyBN6jQTgLmwK7AqoJT4o7NrI8qIVptV2FdsMIMs8besLKX6vtS
WwxIzgyiBeLOqMQOGXzQXEg8DUBfC6cz1H044EsE6HTLpsKHBMhNKsUfpgIiRijAveBpF79FwKBJ
rvZ5kCsERyw+yMQ/PR4oPmVobjucSLgsq8nGbaulpYJiBLU5YmfWvjEJ9CFv95fbXEKuMn2KQibC
6KzmEY5+HRNGLq2cdTu0l4QIPtXxGvV1LV+u0hLlPekzwmGz9wncbYpscqUtCHPHs+U9ihDLAUUi
lz/KONBZ3I+0AHxQfmEzskh5VZKjRoqsC7buHHAzjJDgClSusUkqgZ2xoKk8rhJlgVhLTCJjA1LW
WlcafxLwlXPhPTniq6ULw+vXLAy1QDa+kliNbTMzoyu87sEh2DS5qwZIA2LhgsStQzgtileOHHRg
4YfrPbDPyxv3VRUmGZ35wcGJwH9HdOHqVyXUSRAjjPursg7wRIDHzoSWJrPefSye6u0idazs1VmI
ul4GFNd4YDKTdna0sC/r4EwzCY25J9JTZBnIJzqhxnxIpZatB2Q/k58ro9cLKEh2oUx71m1V3+Xz
QdhIj8c8fx/pez44eHnvKQ7yXDj3Y6Y0CJ3IMIiKlBwouFGq+oXZqV2kERffxiwSZe7wKy8lkdkJ
3rvHBG7kR0BBYZ0KrlIjMy7Bzse75hD+xDxBbPwCjIWxp8xaK50DCG03DmnJroegJLXzsHp+RFyv
qiIjxdJlmhReA7vSPaZ6gZ/8hmTSI1+FQUx+r0upMcF92D/TMIdvedreBR8TVFBktlcziYLLTfRp
AvSqCBlLDkRRBM3gBVrEqiMcYYMPVbPzFCEc7vabwtjVoikW2tKU4Qw4Hwl5Tj1tCSVHWss3rlxq
Y01QyEdzFQrw3XnabXfMbjNha3av2WLEuEWk+aLihpAqS6oOGkFCkXNbeWK7ze6f5v2UydIzy32c
6viLYew6gyH53jerEu8sg0YxmOSJUiRjaQ9LhX0A7pvOhdpdYLjtOiM2jV1MjnMiYVa2iLjCJ92j
018dfwFtWbJCO9aMWxhD4j+FZ85z5Qo7NJpeDstG0ftLZK10jjU7rS6+X2oMPOP1rklFFzrdBCdg
1N3WCI5wGIcpGtENak23XVbjA5QOCr8HBik6ErWzwWlmofeONgrLIWWo/ZwhOFWEsHt8BRHRqbPc
3sxXyhgua90BNdlqEHOf6Pdxk+T37V4ppF+ZjmnES4v3YUMZenLPRnrlNUVe9oGFXp6GmxHQmCBj
/72aVBI5z80tlW8ZfcoZmoMzwUZ09G1SleJh7M03Z/RNrXzN3nPI3GzTgmusGqEJOvq79HIj/d5w
e2YxACT+S2h0HJgwVGjBiOk6DwNJwd+vD62RkCz6SO7CpZ/4PlVFoBlbyDU7sGMYmI7OAuleB2P6
4inlkXUQgOO9E7TJ+L0ZAIPnm+ZiexxHyYOLfjx+EwS/TebwwLrtPBKByhQTa8OdTuF88ZpTh0Xz
IDf8/lJ4Pb+2gw5EfoFMqkxoHbUu4UNqruWvpCwPhg6lk71IqWde2f19h0gMbty2ljngow+w2+ox
EfUHZ3pwUtFoVnIOrNCJSxJ0yiEYHEBo6DNkKNwDW+Hnm8X+G8b4wBMEqQp049Ncv/ezujkuE4Ot
lNs1A5bPlk9SUDyQ2Fy7H+R9Tv3QyafKUpM8yCyfKqESvhVl+vvXiO3TftKEIxCx0Q7uBzkrhA2L
NBc196TpMmyqvp+E/9V02VE6yoJmQp47hq5IqyCqJELaL3mNOpJ74uPllA57upTR52pcpVttzMDH
jRgxgrQ83bUNyik8+X7NGKPreq19aCq7NG8zSicbK3XS8rSRaxUzNKN796qOBbNkuH6wUQx9r5aQ
tj1LT/AgATqPC6EqAB8/Kq9OdSPBNsiLbrGeibKqTx3JBh/VIiMkCXT75kV76ED9pyGjXG4bAzLm
tPfxl0rBPYrmpsvh2/Li8Uoq906rC8Sf/FpUo+uVdN7rjddtBllIWNvb2aEmnWoQhmgFidFFDzqP
S9eHBnbH1unP2DxzjeHrIuIZ7x2zSUj/AGAdVsmSh4bmEALhPG+np3s7yobhOYp9Ol/w7ej8UbA3
9Eul6/5/0uEsTkd/Dqn3QWFGS6sR5J/CFR94OJsD78HdF8Rx0/pLe4iJyRGWRYVQiedBFEPGGog6
BX9AlYH/Zep9kNttc/JDwFqG88Y240VkYiITNIexU6AVDbT6HkzSIUthniyMxn5yTB754b5Cx90n
l9VD7ZGuVOdQLfSTYe53wWLRJMO5w7aKYWYH9QsWTvlpJXpjlttKzl1/i0B9OW2RVnKS/FWKbuV1
w/ioyM88k6DQAGir+NIQ6oVXbWkrPZCP5zbckzvI0ICYJ31KwkKzyCTcuGkExC0Erd3OCbgla2iH
jY5gHrg4bqnKCYCteF0nUAYZ7Ppu1FJVasYvuCB6eSJ4nKV5pf/wcekNIQTRf77NZaHU8E/4xTW0
yEcjhl2LsULWGOzFXc3kx9y17KtV9jgrmEmM3EF/tUpzWadJRiGrt637EvR5XPv17vgtCKNLrgEP
/KYnz18xmGatWdVWykB8yWYGQUiTl/bGdgc9eqILZT1aFUoMfaarendZlhs3tYa9Om9OGSydURuG
OW0GeY5IL+lLCxxgfgHNg9eIwd2UkQaI365qX8Oe/RT/ORnqxoISZRRiRfL48mf1FNCzd7UdWnGj
sp336JQFKEi0n4GzYZy9PmtB/WYfwN7/A2YZCFhMR5rHn8V1BAumxN+Tr2TnigvJPwO3J9LUfNwM
ayuCRMms5wCUCFA+IOpqW94z4747IjEyjaENyTObuXhXaPNdZS16pj+/5EVtDBcSWaeOG2EcTm/3
ejynm+axUtkHte6Sdm+uSR+7ecW7Hw5SPLiqrJ8hszgsozI190jRhvzYfsl7VysfSe5wPICIR+qk
q22jumI1Q1VxQoPhMb+53vgIWzckbDDvDm+jek6ORTOH2DCDK/wz02C7lfoztq/74PLo1eLQ2gqg
njWjkoCe8wMIzlI1M44MmNGCxYrZtuc40RPaQm0WO6eQEqEB/3H7W0uO1g5+DlmptMn5rswZqZdA
LfVma/BXr+MySj9yh9XhH8zg8Lj7FcJkrcDxiPvzqKgWctavL53qTAIDsvmnUD2kpTkGSFKJ1FAj
M5ktTiYCs6xovkrsY0WkczOtue90B0WnJPYjmHmA4FCOtUE7H0outB0bDNyYaBgQaIAWyEx59TUO
naXoogZ8wnRcOHsNHYbN4bzCuPGTerUwZIHxNvi+4xzRIMw1kN2IYkxBNC07H0Hw9ezcKRE/+fG/
H2RqL1i5psTHIs2oGsak1EhaJqmjhjr5Fe4Mk1JBgygL9LhN1AkRgFfliXeQweyt0YxoZ03DltdM
azUqUJE2ZXpXtk8LBSYChQ1it/y2l71sdZZC6/ogDi4ssYJN0mQhuBvn+MVgiSgCWcSynJbD651m
P6vLGs/mOHJzicZsxaEa3PHWDj48mw/JDgdnZqKVSOhU3LUdccVjJVPZeumoQYi0KerIPkZNisVv
LBxX06hmCwQmmZPiv4Y8PD968G5wTKMLkQbiAfLaI+1AsfpoMsueDbhHiTK5JtsaqQeXoXj+cqDW
1g7MSX6pY/lb2XY/jw2TqbRzL1LMYxaY2A7p1urv2SCck8FsZViGFHCRO4K1UE/5HmqFx7tL6ng9
4gEJ1fxn1oEUhhxCl1tbsEKHY4gAN4iV5Q6bnM1Aa6Z5JwTu8yFjGhHblHgsPV5f/1L1ND+liDJA
tzDuUTtcUerTscwgay/rv87CCA0iT6FrPdcbQZdqZ5CO5B4sYo16Q17HtKHJKOv9xKsUVDb52qa6
yBULngfk+QGFPWn48F8zpCCEsUHzjLdcVGE86Mr1cWi775WzfXJaBWHYSBn41n+HfVT36UVc2+4X
U7gQ7hVoDgaMBQcF0ofzYwBEVwy3OvrwQJoVjNht/eS4D+/BealHIuFxheHpeEWjiNcHvjjqxL7q
B3WtPc4Rwp6zkpLA3AKf11LZr3tHtbl2cjvC4rEAUtnbpQDeO+xwSlNUHMUZ0mCCqFnLxT9Q14jD
c5OXaO3w9I1ykTYFCAP8GyUQ7QrHAOr5xLLX2883grWF0/n6an+BvbprqzodqVmWFLyVau1RNEtW
rXFFIAvn2+Ho0VrF7Gtp8ZV7S8JfqVI0nW5ehJKhCABUQiXRA1fA5L5U1nPt2rOQYc4bfd9GL6nw
wvw0scIiyGqBdgmaK4DFDVaQLQepCsIEJk993cGsowwTlQXKE3SpIF8Nu2oMW0BNas3tsSHuaJik
76gZOsoZEgQ/iX49meu5/4hh7a55PJyjC5sTGoIaQsU5rPGC0UV1BaczYtbPdtjo0oEP3mfc88Id
l7HsTMLklIKqLyf6VZyRxVgvCqG7RQJcwUBE/FxOulEMGUTCbY3kwBnvYOQQA07OdAnWiy6EnYMT
xu/g18RsEXOtIkaS7iUhQr0KDH4T08GtTyk8esKV4vAomI48oZqIwwshV/+98Ue+AnESszqZcetQ
NIip+tJhw6fOj9vWOC9vby7pIqqraQsaIcZHV/PekiOgAGnQnDs7mJb5SQEuy/y60xirkOaqzvOf
AK6Fmc9quxAg08t6p9mN7riBlhQAKgcLO+RVadZ8S2UKV7/uMUyRb6SRlBvnCqk9cJlCXdRZRKXO
V07r86l0brav8knrtgvfV+YNCUhfKCFx3aI0IEaHS1J16e95ONtGmmQCOkGldq66oacy5gqIexM4
aFFlQ/h3bOpoTythyZFltWYHB8cAzMp3DWmet/FPH6vrye2Wut25iRMk+Z8FBlrSrkRMgfbNBCDQ
vATQvxmGHBK5iRG7xFdjoinB7PJAkvMrdA5mYqaSpNAaYnNOzOuq1wHtDNWV0+0lFSYamR8SpDqD
f6etWfxHbfeR5MO3NMD2EowEbiYXoDRSZNYdlA9wcP/N0q8nNcsAzci6lDUY6SK5Nr1rfVBNBbqU
ZGFHlaqm4YCwwgUSG4nC4wduuNQwUhEovcrnLyRvoE1kfOKleJgGe1e4daxx5GdptqQAgF+opp+D
tneuiKnziVPrH6FOoFL+jEoauBVs/m8Osx3gw5P9NYz8dBKToT5JWFvYWVZSn/jr+WzM6GVcQS9N
aSpkmm6AJ1ifSQ9rKWyyU1fipy+aX4/j3NVcvtFrlYcfBzCg/Pu/vKDAunWzVm4kBBNSEzgXD6ky
IKPFnCUPg1LelM4/wdAp9ZyGFf8KGlk6dqkLtwyyRxO2OY5P3ENGZP5UXJ6TZ6syUKLXHMiH7sLM
qO38jtDlIevUYAXJhAsxVllPrk6fvGX0RrjOC3P1KKeRV15LXiMZ3tCOvarrc3Y7YEIDR5TuuFIo
W6tp5l1xAYceaHjp1NhHHTva4qL9c2gUlTTL3bP4mDlMtn9ODjVDkU615fOqEosdph3rflzSQ6sC
fUonk59r0HTKwX7dzQmmS9QqsTCyjNEXo8rpW0Mww2Tn55udWFMOppoPsAGqBrcxLdJclzmxNvEf
FivxQV6fV6F5YHpNj8KWYRc7oJyJTNJFrkD6DA6lNH66zgeofcZ6DjpevrNrjgQ8FKQQKeqj6pod
ZOe9MRCLkeninV6OSCtevelFnurYSHTV0gFTbHmOAJZXkk+we3GT1xLuYPTezrPuvO+pecxC78gl
IDQG4lhej2M6jDT8Qg6oocrZGsZHHpQjcwHJNzLQiqQthov9OEBt2u00Pil1FbkI2My3dru0ileE
bfuIkU3RZ2EFF/jp7xkVXsZOdoxGPrHWR4zlqvB5zs7IIrMJKjEY3QQ6c5Hv6OAGyEIfaOfNK5Lz
5zdYATl0UIEKdtaIbPQKkWvHwBwUlMBJ/toujmsIHklFscihOkitdjIlv/jiE4Ynr8UyDqCuD44p
rhLUCodlviqL0KQ7ssZAF0kjYv3LtMlJynGZFxKOoGg1GayZqI8Dz84+P2zYW58iYDk7Q1eEzoQe
bgM4Jjf11Ii+jGr4YF0l69cVU5k8eNLgFkZCf8lbFOccMagdqXdlNofb8MdT1PxXrCEA5KgRPFMD
xyo+a2jJydCLs37CWa0ih/0x7wCvskle9olgsshhk0BSLUBZzfOQMT/yQGJbZ3YOW8gpw0BNJord
KCd5RGMDDCwi6q/xMiu/oNBzu1dYKzas95Hr2sBoBpe+aMo17gsePZldEKGT1XGuSxMY0u9SqrCt
BXADLpBUZhDVI1pSJ1TMRyBkerRsNw8sQtD9xghE+DjZUR2eDbYLT1or6aoMS2kDbggbId034NYX
v+JORmP+WySpdM0/BC1H30F/MRA2Q25Swfd2Kpr9FRmEB2Ih6dvJEVLPsDq5APnblvkkVUBCmLoY
SHtZ5wpNtCyFGodedgqfG6sGBmAfXKr3ghVRRZizREH1L4hY1xnFfQe/D8hxaHpFVo1eK6NXQCZK
JfhITC4QipDz4wWUN+i7oCIwSQno59C4UAiveZvgJfOtsQSEAgk6EPY+Ub6PuNFWLw3GiLFoabNc
OzTudh42UdFdnz1zJSGtlRw4o2TdTl3tVIdwkskJVg2QzvJzIotl6yPc2IEyy2i0v7Wj4oAqC6VS
mymVsIW+BC88lfMFp6I0PKDzDlbNURXFtEadrf1ueZI2Py9jpSF5DmnQQBVzDhl7/D2hpJfpwUEj
4X3y8rTDE3nCdbRkVDjCkKjKfBtllpO1h+HRx0CqNLKtR+t+xUxQObKzinPwNPjKuR7ecIlUqmWH
fH66XaDpOpuNGLpI4mrgdxq6JJMzMrQTZlDaWdKl9tfmWDMYSJ/VaECkOH/u4qSPLhg4+9XCar4h
tJwx0i+5vp5oXnvD6+uKgofm9ikPnm5i1VRsdLcjVfesPtzE6WyQOO1Z4csXfG6zJMpL1p8Fh9GX
VMvmYjO7MCSmAow8YAlAzNqFT7y67dXk9sOCI1UFjA6KbvdMNvin4Utfun5/fKhhe5LsvHn8aGMH
dYJIRyQkfyKUjZZZVBUGWgpgB5GoQ2suomY39SfcM+ngTUzk73gXrLOkd2jjYUge3RIQkrGukVeI
eJX51tkfZoBcKvbyBwSrh3IhYKJ9clBa6IWBezWR+FJjRADAMr7BPKGrxLqjWqxoVAth3Ar+qVee
shs4S72VLE370axXEViE9rfwbomc+KkRTVvjyDO7xS5yfHbtNyYXgSfo3KHhqpWqQ1OuKPD+fWCc
Qyk+9PkYaDvHq+/J5gu0a8OrvFo6OCHWz3avm+O36MTwePUqS3Lag5CgjOmJeIMCsnqDnFK/Yr2r
fgH3eopTY6kk30dwGHmayDN9OTEvNFY/YWmQiCK9+XkzhPuVLe9qBjaN+tXF4okrJZcTYKOosGty
XfLOD65ODa3cREKf66d/smlgFMHNr+kDSZqmWMVvdE0w/N5DsZEEzDTC1vYNVFFYm6L2R3G9AJf3
t00nVLKiSZDtlrVkOrvJEK2cRYXJ4W9aBM9vTtnN8BFMde8UEqioDpyUpo5i3zVbr0ppl3P5wL5r
8rD1S4LonZIZnXFKhCpTll37gNrPqXhkMldmuKoz0Rb0drS1wQs3ELfcNmXh+eDHV2zn+s24e9JQ
0zembclebQpj29J0hrfijzjZ3hNV53J5bLjEsc02n4qVbZjLJUtlwksHPsOQm6YYyFsmU5byhnNs
rWsS79j+/OZGXEQtX9c1sHKjMCAbk/L39J+Bk7ZgqAIdDLLyUkKen4idvpt0+CBhOfp5lOHS2dXi
mQu8X9BzXtAr0kgpSN0+EVJeX01ZQb2oa4k3NY9YO7xjwd77UhhCPgp5lZctiiaZyRfepKAO2Gje
HWbCOTrPpdvFTHfAp/U26dLh0T+BsyG632WjwNUhKNyiYlaZx+uaTLlvLT1JwiXZKPxwmmEZi1k/
L4b2TtHoMNbF8DL/+ADNzHSvR7IXunX8hdRTd9HbJj2WfGJssmRvwZPU/TsSjyb6V3mu05l/4LaI
ijYglu81vMYd5ze29eJSAdGHnea0sdnXS2X2oVQuEaW21UcHmjC8T/auke0ffm61TePHYkRY6kMe
njF2fHtwyz9THZ0AYwwvbhC5oUcX2GO3oEXaJUSEN4zMdfUrEIMmH3goeOvK5JTeq0e1WFYBI1+C
DJQZcDCJxYqAj87VAaY8Z5EC8i8CbbQPTFq/0tkX05vyzQDh49zidlsfX6Q6DdvxetENzSqVSpo+
8fg0/Y9ReQ4TSfSGaAopgx74tS/T9eamnir9+m5Fl/shX4OUVvO7mHJ0fPG5QV4lK0ityv89wXVe
YdWzqPMmD9V/WLRjBWFGK+IxkEeQgLlTAEoHSksxIh9sm99zCKDBeGYhtmUzZoxJ+sZQZGpopwVe
c5QqNV2JONSpMuvoXUtagjgAhNH9AjGeYrFdHQqggpYchPxqY1dpmOiy0wg6fQfyXd9MO+Fsqq9z
6oCMV8eMKZB4oIejKnXfOWkeDQr3JISN/s766NNOx2ziuQrKqDtKyGhhH/fcovVPECf+dk1XstCc
F1K8xqxybhfuwq1oCky822NOXsYJ8bj6SSx/SLqlw0AoLnYn47E9Zi7XBEhfZbf1hNdw8Vx/P8QL
DOdugfU8MqSVYc1h1kSwsCxxAivlJHGzZ0AOZlEKPhEqfla30crrs71gZtJDYmWCCrNHro+PmskF
kZupgocKB+3bBw+Dhx3wQWtXx8Y4Ja2aDwHnuEuKA+eGQ6ffzWNRZALWE+bZQuG9S9MGtfuxgICl
HPytuyF97F4HX17c+YxnZZdp0sZFbSabyeiyAIM601PzxCrLH+v4RtMxicdOJCrQ4V/5KsZPokD6
icfS4miz3Q3+JbaAHM4UMWeSYH0n5FZODNmVzRxjRJWLDiluJy7ZNhoicXmFJeRTQ/2FgJA2ojhB
5OwaItbHxcSZtVew0z6IzXcA4YFOVSrIR69HP54E+Z9vqZnjf1ovv0UGyD+7mreyLf/3b62zglx3
B0t1f93irZ+SsagnlR/sIk90M8ikdc85IP5gu/POThlXH5wsSbNceGG6GZBfGvG4GyxzlB7GBkgJ
11+VzV/myKDgCrUj1dH2plVCfWffbfS5R0dgSWH+ZI1Sue8z23gp59AR4XS2tPf6ERKoKdWP8T9H
qc7YnpD/7ZVM8TIUhP84hOV/Wn0hDytNRAGV1Ei8gbacIS9StRNTuzQJg2/FT35Kz8WBGIu9Z9fI
Hge2I2q7x1B/GGwD1YpdWbf9CwzbkTnyxIho2hb4QGz8hSj8tu6HhC4dky6HWhJ9WTMpWATe8QMy
1kzBDbRQ1J2f1Go0hl/8vpb3NXXA2+7kB8hZeKJadcx2B3pGXlU9pGcau47/mBBFtFygfdt7kD2/
Q0cjofTmBCfHG/pVLAhUf8LJYmOSpBYUDXxTEy/aBYqyCZwHJds1NYx8W0IBrOjwEslfPn1Jjbls
DLmwsWjqbN6JLYaMcd9VxlqWBCUPQdoWIjZUHDOz65qEmYTiCuxb8Jgbj1r/b7AJ6hhk8pP7mTKm
tqXJ9/KJFVApV+uYrzT5T90UkQpVkV0nZOqsp3s/HngcrgHz3sdCh3OE0T9ozbv60//7/cnnHdvC
zg4rdaZ4/QB/SiRKcYPAt6/6qaxv0l8uFJEJ8+F22TRsSZXvzPbu+0eEbLR0d1npLKR6PJ8XVJF3
njpzA57ajQkHaMKvTcH4caTelvHzOvCMAxDtBlQBXH8c5iOHl/+lWVapgnzQW9vbczizHq8a5W6U
mTDYLHSbkYUA2u4+bjYYqE+C++2E4CBQ6UtPJN0jJ9Y3P3Mm5mhnM+pRyjhpFuoN7uRnKvUYjJTj
BalsL/RpzV6j6yeJ0721gY8cz86PeUYho4JjkkZWvkFfi57YC1FJv3ezIvMtleN7/KhQiI5diK2p
ZvSY4p+LjoeUIlZbWiHg8wDrOeZqfLDVmkMCDRGJnk4ka3xCUT3G5Dl3Ss16oN1ueJKKQcPHJFb1
FI2pd0Gk8cu9xWjC+FavgghXLsJZnFZC6Wmm9ZlBGp98f+xTbx7xD+PcxhSwmWZkc3vSgpnkTAeC
S+D0IImaP6K0Ab5ALmK/pFXXL5/ClsI0+rtjDJQixWn4kFj6LKf+SQDvSEw8C3bskjKw6x5XnhF7
gnQmr0giwIHFLK/ecM1RIIWCG3yDIDZEAy5WVLCzzT53i3dY0TZazZHFgJnLIMBMXyoY42lH8xZ5
qgIMuMA8aiVVPITpODKVUysKqtJ2ywIpQBmKeyRqjqAsQcmG5FVE6/adR/CzwVI0BOT2J5lgCNkH
sMMRVPy0Dm0ok2MvVK4JwpLPMYy3qK+zU7XLao7fYf6K5+wEEXuZnws0NhNiC2YYBrspMhAUsiYe
dlElIkPE6kejc3ctNZTHpxgvP9VAcHqIDhG5hLOYbRViPsZNbFAV8+iPuvF8qSM6orYGe+4XVK7F
lNSt+UIIyObdpS6bHXAqWR1/ritdBMWmVAUi14v/gtSHSsZykG1pICUhLdD5NE6X+n4jpBJfKhI3
UOgUV1hhENGzsCpGtScT6wbHlg091q2E8fPmL2jtBRW7qWJGqKSuaCzOBvT5K9D/gK8rL8S2j44v
PepLWZCEzq28uSv/C4GKbLrLm8mM4tbnVEbT8RtaxGgihHeN1pcEWsf8SEWPD4UuG0KfeU9Pu9L+
pqhnOb6a1hIvWjqhbDpI6CaK8kEyD2KKIu80YyTaxzcD96YnileDdrbOcX+qqjtWHjxkqT0hpv2c
+53IVXykrSwF1yEQAYw6x6D0e/6/JWH4bi/LsBhLv2rpa0lLNxq+VDbZb1ILD2q1J+QxUnbbD6wq
0aast8p3+NACiA6nl9JvcRXxUDNlPsaLPcMW4XYbblRaJzh92yfJcfL6JlcQgVGgcZP73bAI8APQ
Lz2gPmGpSZan8e3hUKnS0iFOy1qs3N3FWkNL8ca2rCXxj4PDdBHbOpQkBN9pHDYPlLqzVqrFawlF
vB7Yv8zk8jFO7qdlGZXGwq+oH8vSC1uFeFrUlv64suvIICE5oO3Z51Lh9DeHXMUOfB2wy4p8K7wu
w9we1P0wFox43c3QaDH2rcxnSmtLZR3JU5v87B1HMi6M29ke6G5vF5Ozu58waKz1xFPmoPDxJj0c
7ay7Qn6ijnxI2aZDi6jyW9HExYNaoh4KvZfl9T9jhdfFBHx9v07D3UE4lGFcLjLhMXoWeBhU7YD5
9lPC9GfHdOPk+3XSnU2IL6X3dM5XW6rTeFZzht/b1RmCJxptTy0CZvRRk0y4BBmQtd5T7qrmJz1d
O52DUpjtI4KQ/6HPiL0VqXEn4YI8otMoa/NM14E1EGKD9Zc+QLl1PVS4H+6NllhM5vARo4e0FfUI
zo/rK1RtUNx9LUfHnjeNUql+WeAcs3epYRRAEch4vxsjOm1xGMlrkSgYd7QEmntfp6oS+STsNxF+
5DudvKuq6GelTOW3K5mweEELrksPkOGMHzl/unC+2tVPI6yLVHOxiFMUILuxBReQ02gaNuRorb6T
BbG8JoINtlM3FMJam9tm7Zy9omXPjzsGEpOSkaB07lQRPjTooHBwrrwe8XtBglFbSkVtAO4zH5t/
AGCTZLa0RFU2dIwaDVTXiLi7p4XyV3MxEyek3Mn5o5Sl81LWLPQXJ1Lo9/GSHf2u5qeeu4zvnGLP
nfM7lPJzegoBGf5bnIci+vMLR/57NDD8NhDWe+lQjnOEQ9o/tr4XrHMB+Cu6D3had0jiWnDAdr8u
rElJ3ogcthJBryTaexRAiHndWyaHt5YHSrwebnGh/MbhXOf1SZfzeQaIeCjGKXycN6EW2/E8dXvi
cGTI3nlYA2AW6RWymNClDiu6dDrWNqz8ipuu/bkX2MDwxsBx/mYM+DqJlGKGsFwArMW4gNz5u5Tj
qmHK3eNyvfkaBvRa3yS6bGM0MQb/VpBHW2MoosxT9NMHhVXYb49tlqOiQL8DSozdSQATMiqjA0We
K8aPNSva8wGFHVjCYmTNfhHa6CEXOid+9LauGYCrHdYpV7q9bnGDh3qi7fqksOexhWOwOU3UHUY7
zyWQ7YAcVDcqwDFufxCpPY2nwrGLV6sHo62nVUPH+OdaRVVPbJHzKiXIFmSBy5lrViGxeGNB9q+i
HZEHMRuHdBJ9ho9j8akF2GvKvBd2Ex/2TsdEQU4ivD4mPY6MYcmzO+Z60bVKMcBgsgnNGqoW9iUp
smKHYAWCbensVepEAqCydnUL/8sdc1wgSr86vxPBMitrW0flrkP+Yai/JU+EfnN9FUxDRIvVSdvw
sxIt4FzKD6knwVR7IEsgSOTuNvAkv/j2N/4d25qnUyAGS8bLOJrvHuyoeI6D1m0b6MRmysAMlcdo
8oqzskctXHDqFIcXFPjPCJNdlSC0vk57SqygXiZOs9htWEkBOfy9QVZClvtsWQ+hUFZC097/ukAT
zoLkk2W7/KdSRbWnh24YUgBR6nEIBEunqa6z54GAtRmWIBKu9WjDVlhGXwbpZaTzT2mIjylYGLFS
l7/+iDZuVoDZkkBkCTd7TX6QuBro5AmxIDmrTdE+WrHJlDYJy6a9mUn0fa2f2nl5934Kh0nIWNFn
sQTfFPw1L4NDFftbVrUpXE83njyglFZnbs+DH7gC5slfZB9IINf78Dlxe4uxZIZ607+6KUBXQlPj
dse3D0GQh2EKl1V3WLUaBHRgqfN6rxLCLxhnQN/Ph8yVU71S6NBiKd4fZri1/j6WOnmxQ6KHrhGi
hxa2/Sgf5YOXYCaclqOGFRAPXWeigGej1FJME+9qvWyuxNbLOxvloSQmV8OSwATveUlnJKUATsc9
N6WJkQ/XV0E97xhoTuePCdFGlH339W06VK7TkMqphAt23y9NZIYQPNJmNc8sh7t11u4T/cEiqtDD
vyvLGNYwjkWDnbGO02A7jzZ5+Fl7wmm0kk5xMuv67WAc35MhHWkYjAdaqnC91iRuq/I5XLLz8NcK
fR+7lk+EkPMoG+bu7JOabn/i9W7gLWS3TVBmbx9puIh8Kw1tGVISrYzvd3verEHiXvgKhurkKIvY
npjxYv9pCOePqlE+Vz+q2Eow/btd2aDqI/uoGKsx0pnfSCglJM52PDHM5pwcfIOAteHlobg1Vo7V
ot7Y6WkoNpFipQaSrget3dEokFe+vj6g5xdt+uZREHLRij+HDdOn4enqTZHzEhlinN5yZX4W7gjA
C3ym3rkaDYs+YpMZ0lSrt/G7M3EjzAfbJKfy+GKqh8MMlS8hxX6CMn8E/2PTmHpNDfB93l2OqB+t
Sef/qwFmpy2ugDXsMbeYYPpNg/LSkhWcUJBP/Wi+U5avvW5C6f1rAcVmXIZ3w9PbkacnulxFEO1b
rG7QfKjqN3oHdEcSoFRWYsabIZKAJnv+EjfQtdc17NC5mwNsIobL/i61wzYv5yRLGKldmxci1rti
7nmPU3sdgwSDHgn2Y0PX4zCXC8qwaUgjymqrYa3lm11e2h6mrlea4dZk9GLzxJ1I5wAyGM4aTRTY
RLmlEO4SLMyNd2sOXnh2AcbqZJPbZGn6MupgR2f1bYT2J9a2z1JMOwo5PNn8dOmda+XktnFkoX13
xvpwH8M3jpRSTUJqZpPRmYCN1aTysRG6h59vtPOMoLhOsZ0/BOhmg8gAYlM69gQvPga0HiSIUDnU
2AagRyWZM2stzWSFiz8RCZyNdHcTivlZhSy/toxnE4Av6hBQZ9IA40UrkofeXYZExc/w8JC3+VSh
S6SX5PkZlOgw19lc5qWjcpmFWA7Gh6WpyumDHmLqiMTfz9kd8z2QyTmMZfEAOamvXG9vsNm8DEqb
m1C7e8zQ9vxD7/g15WpMjlJLuQZc42oOHfkxlKpIiUBquNxUL3uEXlIE4GXZRtzfiSAt8PvtJsyz
3Byrxj+eei/TYCA3rBxG+agIx8I3v9REimQbT3ioVCk01DTHzRAKf7knICUAloLiB1kDshsZjm+V
30WQ2fOwl0FHApsaHZySpITMVG5yg6rsuuwS3xg+2SNsfUNbXdm5u5jAJEqm8HZ6iwtnNnPGFf+y
6zbcQyN6XD6dVtI0ImwmkslnxK4h7Z8Qa3Ui18h4KHVcEAXWFEO0/aTuOA76BGgUxLZmaNvU2JJc
QSGVIt+S6+tMKqg1Ns5q8VEL8f3nZ5hueuzMa699AtTDdmiY6E5Cx3y9W36TfXreGruACdVCl48I
ROS+8LqCMkGcwSB9x3hxnnQX4OcH1iFZ7HDi2M4up8ThWWy3WeA8zW2TXmZSIF/aVPukVw00VWdM
gyVhDc0yhJdNcfDJYS4rd0ug6OBV+3SlHRTGbpKeD5JYApG1AmNpBV3QTaxpX29qR7CioiJAFX1V
dolrBqBKImyu2Oe5QJ3OGFgfojt/ET+R/EpcYWvAlXxM3Y480AIDKeidSB36yg2Q6hcbgorIdmuD
tQljs6vCxB30sWf2SkaHP1FPD4v2WWx6L+vBo1twW50btqLR8KGXSWKbsC2VMfQTJEIYynUfYopI
jw+42V5sJbMfBwZQ77poEmgGbtf8XC63z8Scgft6YSPCuNIeOJ3pVQVWt73y9f5RlMo1UHdf1F/7
4WwGsKPXe+9jLBS8ynDKCHBUtnbJvToDLrNRBCm+Ohv0+uW732nL+YyAVyxJcs+lEeoIO4XOwjBT
xJIhd0RzC0ykv4r355N4q1SgICN1ybkFwCKYIVdorz6X42Kt717fQQ17KfDLOCwiJgXJL6f5WIzD
VDbDntfbeZsOHf0lRPMF8AuZxqanE2t0/ZzOLMQDjHUkNmK83HS98DnMAnwYcfjHHdLOcNuZx2/n
QLZ4OnzlMt9YtemrIQk+4bmUHq87nB8Grqmqrse0v+Oc0+4dKn9D+bR2hYQj2zFMyCmJ20UXa9YL
PI8PeLYvR1lhONL/CkrdY65/TrdeWFUJobS3DSxciDceUPoRQqaphYILII4PvT0sEQboTTOV0s/B
iZ86QtD+gnU8m2yQpQktA6Ln66fI1MY3dEUwIHK9n98G/99Asa35wKEJNF/r21AXlYTPxecg9N/B
G31g/Jk6OjRs8fyJBBvX5N3v7xmVw6HJeHVhHfQ0DsJcWc7Ij64lmD2K3BKx6mV3OR9ST0eG2vE4
KYncmu3uZsXrJdXt1miKzJtoxdbMk3EzHTAGHaJZFbAyiwTeHGWfsdZMDuZVpSZFfAHPDxVmvOnG
1r2KUp3TgBdCHvjLrCmGuAiGP0qjB/L9Z8hJHsBJBp5rrc5c24QRowX9sLjahEcg/OwB4VuLnOO1
vak5/0fY9tck0ior0Zb2cSjapYqmHQYbjvdYYBTTV1dL3tQo3I1XOQ8SNJ3Bwa+XNbJptMh7W1Q5
arw5+qJ0+5t352Bfe67rE+08lJkT7ARxcbRuwe0bh3z9CGPzWnxdLZZkMsLmgsS0M5ReFEZ1g6R5
R8gfFwAktbpxpp6iJwYa+MM3yEA9Of2bxjpFrxjOkGu4O7FB0kz7iO9HY2tEkmBc6hcAv3o2WnLe
qoyJndObNGzyiMrMNaoUCEP0SNXSZB8TyGXcN7j8iLv9zdcnyUoBOn6ihiH6wdSILX2IQlNmKY6V
vBeWyhDdD6OPhv/8HTpKeAt5ow9x6rs26QBUEyXOU8rTkMtbBMmE4D4ZoeTzji94Gm3PvcIJkd4Y
lmbATBfTw9g3W31NzsYzPTJ85QfyjR8ttmsgUf78gA7gyAH363wDe41AMEsF50QfO3k5WY1ALOeV
QubGDqsvUhgqtzIrVQApZZ24EfTaaQUvzv+GJmheU4NvMI0DqC+XfgohwdMtrN5YsA1g8oIbYNZ8
NNhX08x8qBa1P9iielZkBQ/+aVzfoaFzkixN6TcLzDpLpSFN2MGmGLWCaKRe83Tuppsen9Gzqgbk
Ggo9+/Lp0YkDaI3kexwyKci9Z5Ns/fAsvCrxIK4/U2ErDQzfNo+JtjniilgWb/wZbWLVAosbNBaE
IHdkgZ3EfRFbHwB8Z1o3yFYP5clV+gKJCr6vTbQRB042LZT/MLqGGMgfbPswwxjVAtqsnYHb3LIB
ogQJbGyCeNdnK6vixoZgtt29xGLnFqm7JL3OhSLoHc0Jnk6rZzC5fXdzOVTcgLd8K6wcKWkh2jxX
h03KxSgF+8xoaO0Im0wFgoC4gF6Hqhv4f8NSK+vpGDp6B+VilTb43nWrAgpQ1cPzggiRZHbDi6Dl
JZVnpRudlN5RsFOPcVAoHwt4GTl0TJM7BnwnkBGSd3E76zGhh64d9XiYn2U7/YGFkqbZCze4edSe
DDHAF+UN+LVabFsIjeUNGR3G+7eB9iuXdA8BpqGX0KwkeF5QqLdxgfthC79UMAwFMXiXB7mYZCzD
86L2QVkWunNwOwUGuaMkcSNmbIImifRePpw73hu7IvsXr2PkrxYqtiP/j5al7rMjYDPJQARdZKbu
pm0Hc254b9kBJDKab6SnKPxcMCVbCDeOKpdhUVLJV3dWvcFpFLALBR8oFQkgdHNzp8VRHsjv9Fsw
0Df6MLicgFetsu1H9+r0PlDGx8HSMpjf+xWbvns0wMMBMQ6ok+DuXlkT9+j7keomDFgjH8yuGKv4
AhlIZcQaEkIJ48Ap3H8ktQfd/YRhNxQhugGtzPI+1QDFlK5Gryg2WKWAh99axb3FCorgLpz6bGR1
/cWDtqChmiMd5XHkretjBD8R45ESDplFnP5RBUSJwUCPPK+/hHUPeoYSm18MJCtEQelFAYkDtFTv
Zlc0JMI+a821ZKsHxdaKzhojBLOJZGQMqXFo2ifkBtOAjgWn2A1Rm61QX1aN/tiGEVAJBDbp3mhM
DfxWKZ1yVFl6lzghCBvqdSMXi8vc3BMX+N+/hn1EUNLDv2TQgbwnq15E+w29kM4VG8+WspKr7ZpV
uKRc4tSVbDsGlAq51dDzYQvPShVQL0gxRtrSnVSWD/oite4U1HA9VERLJLQSmyouRwtVo1zppMPK
VbRZUDoYMoLMmTuTr17CKWpx8vkId04OVA1zP/rKd3bQYpXdTX7nthdDT8tQjFXqqEeStjR7lAVm
cz8SizLF6C/vmpQUfJkuxFuSrDeZV+X/XpuZM9kEtoRt5v/G+OKDJaKyQBc/hQnma1m5XYbwvz+Q
3BSXeOkTPqAklt6THhL8lsj0UZeGwvRvJsCUARC81EByg2SeRVFI2twsTk1Ascb8FtautU0QRUw7
JgWttZHlO4GwvMB3za+uMWa2nZAtQ2zIkTtlcGurXM7EYRxCPdXWtjx0uxiu4+ZUzkvrjcUv3nDk
z+MPauAgM6Am5v2KZo06F9ThxMWC+8oApimNMJSqsQ1C7M2mnLSlzQd0bh5OHE+e0/gwi7KTNEAx
leL9I0BCcJ4y1KCwjBaeLZdyF32tI/xHAYyZYL7r2OA2mcOuX1cqL4Zy/g5lNvNqgwwn9/LpwJoF
tTQf0HdttubWdXJyx74hDN3KsmZ/d6CYeb4h1dK7Ow4g679BBB8wt3y+RNX/aLBvA9+yXW1ulvQX
map9bpyjcgAXkzYYRCDXDJo/K2AhhKonYJihgnvb0KGpCUsSS6CgW+4U+B7pfK58sRDr+gnGf5Os
eYqBUWBlIaLNuviUHXutRkwMehBRqjsYwxASswRttabKhxhFKfFGEsooRvWRPwX4Wve5UEYKt0WN
kPKFxc5jnr7n3l25aYiyv59hvhUvBHFauQ71N9WVcJ6MOYTLjtUkKxKd2Mphgb6lkdVVM3+Uc56T
ydujCCXQAodNfWZ1V3QJqQ4Jpfo8EDcGDgkp4iNGJRqTiXcPjbx98cZ6UEBjaKlK2N9H7WIW8Fqz
3rJKmMPF6/rZg3mvDU/rpxOBRT4Wl1uJRAZIkqVTRydAv69c7A+8/lzh5Uf6tTZDazJA0h5PiUlV
Pp1w/NW+3zsPdsaLSJCs5cNpFLqsbDuVFnhFwc57ZT06MB3U+H22LPSYN3g+g9ViHSsuisPezmOq
KmQk+U5ulYxnTS9sbkoD8Li+L5Mv/fQhXe7Fwh8yqXnigyEmlMNeB77g9ZiMvpg0eabNS5BzEQp+
H5G4myHcDfDW9vpOonyK6Jb0Bvoy6YWTHVLYwfdoVVrXtqwsHTA7cLqQizjv+sAwto2SZIvQQN2I
Fy0GqLrMt+ZIj+v+ZGv/RayGeXe42RZhfUM8N2BzchF9Ra2m5avxHtp26Fflghb99oxiAoyjb29T
+C5SHXcwSQL9Xz7I3jHiDPbb1psKUvglFBhdiQFy2AskdQPwObJfSU831XqM/wabypm6ClJ50Pl4
WAv8wh/EGo3JY+hOQ2VUj7A4ENehrBgtABRbji+ob/Y1klavzgdlZp8In5zVTty47WXvtw/HK1NN
WU/tV886CcPCOUs4rCZWzAJzkZOxujQRCR/C+6uu9TIVND576IkPcYshVph7xf9xXYqiQ2CuONah
sREMcaqPTHciwqYl6qfbA60uHLzwNqhUoKbJbEcGnfCQ4qHBbT46lc0CXicfDaqCg+vOklQW2IQH
WZpB2T50Eg5kAobEQgRdUOJGOLgmTBCTNdc7Dkt0xUXeeQPWDtXVFGX7EwdK/YWasx/311tYTdCE
Tqs7WPT9RvwERbrjEJ6Dj/6jlkwQu8JLnkMghmnrO8Zhi+R9R0PObvW5WRqqBRA8aGsThD2+PacW
JvWUrt5n1dd+IQiTfdx5KcGg/AMXEJYmCNspyuxb1XzbaCqUREDcrk8WHrHBTuArPxw7oTGFUqG/
5u81EsdN1jUxpsNsAauEHSh0ntWAbtkH+DU28WhMV3Mcv/mroaZV1+8hPjMtj30TwFhv+RF4e5NL
wf5j6mgLrjNwwEsAOA+Fm7rLLCysD1whdvpxp84Zoug71uXLUKCjZDv4hrDfgnBHYwRlnl+C0EcC
WXPSv8v0yXtejfM40f8pAbfEg35fkrB1+ZsGDp6I/f6u2Cb3cn0ykNGQJ5xfFii5VTRfHW4f7Ue/
QUzEFzR32c4ZSRmLpFVM1j4QRwMpw8NI257SlvKOyNBRTMc+htFFuXJHmrAquUnqMmQ3jq1g68dh
NKWi4n3ED5f3ZF3Vdjr4Vnsk0lIp0d+OB2srvLZbftrjA+B3bHvkfCOJ5MP/tiRcBr+Kyg8mTNuh
VbS116hfvXvbu7AyIjfSYVM2vqp42ZX4mhMVnE0VWRF1pCeGT5C3cEj0LGKZqcjjGA89i/Dp/Xg3
8GAzjLoEPR5Mxc1pdeXvu4WMzBg8UWcmkFa2wz/KiJL4geDL5nTf82LvtF4fpOMlBDshz6U1JI5t
XUCOMl0FPieLO2U3Gwc/QzT/xQQbo1G7E+FSPGMSwrKh5Ny7Dshr12+z65hd2nz/nuni46Ep65BZ
aUbBpojaLPPILeKbbOdLXXMufNW0hTqnWqZS+31Wm8W6uf04c3oVUdoPFeWnfwCPc9W2wVhHdyhA
/kK/8xyVrttHPHBmv9I/mmcJZI85s3yAmFeWjuDDbIAbxU6MpmA/lC0lbkeO3YT6aGMRRuCLJF6q
IoxrWAWL6GysCwS449Jw3NPffwUKcbtQG3SupplGLI6HZf5TTTLcysRIHN7iT7wRU/xQM4WedlsC
wAhEcPcAniFLhZfisAEdnswNwCAetwhhavD+Cp/Cw1l1ycHLs12b8Xx2PGmGKIsmT9rs7bd1Cxwv
0yXngyssv/PBSMQ7zLY4a6xcOemk/Eon63O0vuNQS/SIPQqcIutTDMIXsE4RAKoa6MzbeWiUJmy+
R7Ol4VpUwz1mwKz2+yFb1RtD8ChxmLopt+soH8Dt5iKoEzdvTTbD2gsjDIy6MOYzgCxl4RahobD7
7HiHisg+Kg1un1oSrU4YZ873BEuEbYo/ii5mEo5jjIEACEOLRPtj10Mx1J7Ed7mDrJYhvSjaH5nb
F5uYUgMNAwSTGUrr8rRIv8z98DetctDkN9rGCG9MeqfDrPfp3khujjA1LKjrAJGLT/RKPWyJy1IV
ysr+df3VaIJOpkA/3N8ODbTgiz4O/RTx1ao3a4cZUl6KZ8ePM3apRLI7nFiqQS5LX8wE1ZF/ygyQ
jVBoVQzgWrJq52f2E5WveIAIvYIljbD8J8LyHqGgLVNRM5E9LM5CauJVwOPE0asYAuL5wVpEAWua
2K4ho+OWwuXGn2hTVWwLAtkDZ93ug502GvhKSPHHywcfjHhkEpi9WEs0NQkUJ8uqc/oyHX42M2Ry
t6jp0fgOEDsf5lLFY04UuKVZDRl4mkOsj9MGBiJMD3sKedokqnRc/nR9xcw75+J6xHN+AqIoWJiH
oDitfix+J77mMV6AKZZWqyNOC+ZZk6eidA5nZz7Gk2a/uZPmQ2vGetC9WjxZM5CnWNuf3/umYcMV
ws2jxkW3D5SBvvscwVf6/WyHzYizX3gbzVYnIQBrzrBQxXRiRHDoMPYXvGCUxaPtW4VqdJ66DX67
X0Qra/0ApW/ETujmd7p46iUu//t0XTYJjxANNbiGMpQwXpnReuIYmO+rPekD3034fFLL5Y8VDHjA
d6tCVCgPCOaCWwdfFuC+iHdIhCKLwu3I12q18ZtkvCn4syXrjnJQi7Vzke0H7J75erJCFoaNjlK9
ZOV76h+i0tWMOZST6L8WAAVovUfdHoFr0Z7I1iuYOauPOHHo495ZU0fT6ZicuTrEG9J7/orOdSu8
9OGFTObA2p6HuB4R2V5zCIop/KyMQMVfyWR1ZMvsfat6L/6IGNY5cW1SCxc4/Yz22nTMyn+nICqX
EBXmeFItV69b2V+epsZu3JruhtPAsaa3F9TT6M1OuPTJGOS2+sLl/eECObMBo+C39Zneoz/YfsL3
2jeKMfZyC7BG7XCoyyUve2YM2EVPUpc9KuD2yBx442pF68G+mkvY7yyqQ/FJkhDj79/X1Kql2spD
IzBV+7y1Xto1prYOYkNq0PtIgmc2aveFAVRN0dEnykofBO7Yb9/hxfV3qxOSLaVDr5ZhEaRy9XKL
JPFuBPWHFzxPnCAhJbdCocbpJzTzwNwGxW2WQmCkj6i7OqCG+w+ccAx7Sfkp/ffwqmSBK3fTQhi8
asbtHlJSrtAh6v8PiPDnJCfB/ZIWjRnq8QB1bi/GfGIO1E1F/wMYDMiLSqbZg4f6uI9SKlD2E1Z4
+A5nCdAgWvVzqVv+wNUkFGWk+k3G+C5keuhkC8dEdXGyejrAkQtLaLIEInHVGSvH474suJd3sDKu
JRt4d3JyH4W5XbdEow8Xt+RqdZW5kgySFkBRWgPJnQm4NZM0MGnZE+TamBBAuVA+NcErSCkhy5vA
8Zb0SuHU5OYez36soxlmXisNVd3i35AbpOW7zqKSEJTwPa6axkpXcc+a3BEPBFEJpW5QJsBekJx/
fODEe/Cu4Ha2noFvoHSnNgd45vNO2wBiS8PVNftIPkHZ+wBcRYpchdpaSF0lGc9r1b6PlYwKK90L
DeKq+zpN3nRA+R3KLLILqXqd8BvyiYHcDksAvdkiwsfwSHkwcDNN9DdTaR3gtf0/k4WVklLLrbef
W5ue8zJbmPiwT1S2BYWNKix0bPJ1DtyCgOnugCkNsK2FSGHL4VBNTrjBos/rtuv1h0kwFcdphNul
3j8lU3uFWNxoS5HT9oi7FCfx9SUxZ6EIjePi5FZ4s4Bpukv+Ejkoyk6vCTQSz9+8EjvNySk66Y7u
s+rEWgdWFqyxwtqkZeP6wf+S4lCkxcIWrbvV5SgoCkEvpPvbdx2OGqr+2I8zHSdqmhRkKn0Hkmlc
M9HsWvXkek4qWBdK4bAvO2+mge+aAxSFiHMELHMNJQ5hA5Xxsv4viViGSxzgEOZT0cprnTsXwbYm
ybgV+Cv0rBHfR0tZOi0vwkwahFahVKf51yssWs6NRvSomfU7lbkiZrib8qUiKuQXVMSCTxsdmsa+
fm4l+1Ko/R7FYHkdl6kbbfWmH5jeBcfFHGeVekk1GUZQJLfb9mkg16w6GBf6mYUmcvOkFwFSysb3
UqtHLy+lJKRMEb6UL2O+JqtQS/v8kTTgalMxEv2RWmZy53XNKHtr3v/tCz9T4wpwO7Yc7AolcAXh
LvRQbAFLJkuW2kN1NIDvHTVUp8f+phjYsGYBALlqP4TTI0yzNmWBY5SIwhQyfx179medeBt/MGr0
2G1Keie5+UWiawgtaGwe/uhsJdfZnsmkJobGQxeqWQddEZ0s8s6SEQeHz+XazV78v+yWWO2LdtwF
9GiLbDiezvwTecQWJpgqqFoohVxoCK8o3QgO/WIy1Ksd2ynv7+1vAneYZny8qkmhpzquJm7o5OUK
IG2un55XrMty52KncFyYIVILcnsWSg2gAoDPhXgpetFg8JmWpwrbYxsrZ4IY4J+tA7sMS2MGoov6
4AamJv30mhRLDEj7w8Mqnn/P8e6dUoB4//6Mf7uM49P5Rp1dCGyT8C7x8FGn2Y8HiCD/KT2Z9I2y
UoOxGomqMcMU67dQoaSwdXWUCGF6v7VVAkbQSgCdjUdW51DViJLqBGWJC/4OZcqyv8CkchO83ItF
J3cUuwqCEqSUQD3Xa0qvuCMfAuKjlC550eIJtsIl4afyC1P7aFv9RuuEE87ePnjB5qyN7CsNbcjq
UIL8xNgN0iLtglHQyjdo6dDayV8KhDkhbKeCBzJZS2fdL8hVlqyEkJL0wOpeDDsfvnT7QM2B142O
9jIgkfvl/z6a3JRdAFG1u4Xcmybk/xm3SUSPqId+bfC80a1O/Iz5dCRxMpTIt7dfrg9/LZviY/f4
JMthYO6NZ6zgQAUWHVI4bFKxi9Qr7HSwyOgAfNlToh8WV1ulkAiSOzvtF6BynTqkajN/+AgkaGod
eB5UVSSlOYCPQsqyGzS+WGZf9FFyxu8DRufiVNyfjcJ4vzXPNYO/CuREyLzvBUvO7uol5ZptyrFC
TBIROjhIDnUqKriW/EdQ1G6hbdk+WxVD2nzk59rUlWfBux87ATYU6ut57EzKU6Zu+FZ5VinHWg/f
O/Hy73k0e+m521/YYO2+8o9ONypcnDdPNqXvQya5qyf93qwUcnY6infghRKWEn8ZeQSgJO1/Po9V
hWntcBvCc5M8Y3pXjc8QubImu1yZvcBwtNbqdkSIfxJnFNGMOZxL5wlniZT3ovB08b/JoThkm7wr
BTCh05RK3/tS3L5A1uYt4oQ1ljwt9ltEv6oyfO9dlr/LR6uBy0Tp7avA5lOUUCX7367UOkJdGFl9
o9HI+CpcZvgRLKmYAR+StJH3Q4P63+D5uQl9DyclLoastJI7vlVSXPYtsdaA+79JWJOoNBqeVS/f
DP30+JpCczOL54i+GWidAEkLoQLh/e/LG9w5dJNcPd9qAE0CVOnGe7bWxaiWYolHZ4uku0lPm74Y
MfcqBr5rG+O1tq7JxlDKPc8mfH5Q+ivVBf48+wBIxsp1mBWJHSeIEe97otqeszssz5VusLRcoY1w
vZHHHp4gVfotPoFfGvbOv7vzLe/1+HhfaM3OPNol+LU+yQ3yqDsD32tY2lk+cPhUaDS6QEkOsp4r
RcLR67g1m2kHrQLCQQOe44cjFkZREwdKEg8X93/BCbb4nO/xhZnXBDKVWqNphwudG8q/vr3z0Pph
lECLOWnHHsGRfY2n4BQqyZ1NHLKEJULwsIcMbTmeIg+4rE5v2DawManIBShw7chzhWU1i3F0Zprq
i1eEsWjz/3U1kD+jMpXN4DRZGECx2nU+c61XJHeZIXFrupymU0DPI02SmLKEgzpRiMY0vD1oIGi6
JyAxe+V+eniNSj668XSQ6LxztgAj7kqm/yJUoZlP93fvBrlRD4pW/vkvcLkZv1D+HHLIGktdZdAw
ovaB2cUoPg0Z+nr3biIFXUuv+cd2zWtEL4X/+AYIfMNrKZJkFkQmFsFXfvDqpUTcT4NpjomD+upB
CmKDdbWGombRW3hM94TF76FjCoVD+KFqbTDrW0wefwLymtbJh003Cih5rQStmmG1GrsiwwjIIW8L
NoWQFjH3lKqDthlzNeCvbG1+dQipJOMJicKF6pWIha83ypJma81kGqWMgiydCn1StxbKaY/sRwe9
GYZQ53W7S9vnnWjZZc39SRD+JJ1RCGeARTorSvgzkmUX+o6J/79zhEHvVRGln80xixzf+VCjY5WJ
FrUplSqw/Ey8TWFqbupvW0xlAii6jq/O+OYmSnW1/T8TC7jeujD64PK/8Dr2QSJ2dpLZJXfRC/AW
PsJScT3ej6LMnungicDAZMYnX/xWayKnA8FPBf6H5RAxlKFmWJlMhrutodBlTgs5KjOzRnDEmkew
82jZMW4l9m0PYlXMlPG3sQqa5xrQsl/dDxPtKYUwRDj51Biw9lHkt51p5IZll2+JBU+12APqdAyD
NY3Nk7DA5erBEAg7EwIULDsTFapneunGttric9MiEFAYN0snSYr1GCnGXW31VY9gsrv+ebCHEFwf
MmD6EmCeBykRQ89vhm90eble46IqvkCirF8yB9Hts3ZrlIE6adMK9S6Xf0boJcpLxBE6iUeg4pOX
s91rULpMfO7/MZUw9+LVGz9z3e2yavRye1k/8/pqtX2h4SIQKJX5+4JQhoJZWLaGAsShG/PR1CGS
9Q7CgXJ8V+jClagU9k9EpDqCzsm8et8tdq0an/6a/1fgKh8qXPQsUF9ZCv1/2I3ElEKuQMlTnjT9
Re+0ALOOwGgEGr7KPgyVJBRbt+AVDF3octOXT7xgmr7b3tOXYUj7Nu+5M4aSJELfev1YIhF0lMqS
c7sc+BqdgotC55e51AFMroemz7cLBL/5ADr58kDYATNTPy2Y1fjLs/Wy0KQ4rHnLwE2NEqE9m99K
xHkwlCFf21/quDIqOaiRPkhjdmip+Qe6Q6GfuVjlndijJKfYOzXsCmR7qfSMzIQFHzdChljrkSGq
048Di+ZAWZJ6F8EIBLZn7WoMgdEVXJewnmt5+OyBKkKjlQ9xESNVB4IkpKY6xMtHkbf5MvJiJiGx
YNsNEyQmKt7JPhlwVlQ9zlXnmE/CW5hmc8zHdse6pAO8jHXk0oqJT7K7QJMpCS4MAr6Y4uCwLclm
/CDrRinxq0KtII+nCwZOQjD0QVPEH+LHf3bSzJOAIh77GBHviuU+SzKcR/ls4TdClgtq7/IjVmrl
/iJ3SrRd1RCoi0VJIm24UlzDoH+Bz9caeqaFJig67Ix+ju1wY7yzsh64sWaLUcYhrsqx0tdi8Be1
rKMeNqLj7lDWdlrRHDsLEgs26A8+Kl1987iepOKI60M5zlS9gj8epXlR4lDoTdiuGw6aMbjS7uVb
twlcVoYGt4qLlAQjCiPchdlDVFl9dNpun3HYjg3mXcQI9gK3DzuV+6vtFJNoO9dkiaca1pgdRWpc
Dq+9VzT9MzwoZ+FlkRmTKChsxZADMRu47/UUcmgimwj29KoFsiGmOXbEE3iRT44++U+6r0kaWvo+
NiwNwLyf+xCh0+TRoDOIIfNmS1GEGuLqWTO5dvf27AJhQNDmU4ISYVHppAxTbS+gMlJ70t70ngcP
YGIJmyp2MmZ7ac2C+iKkh12yONiM2UXBwFwU5CAoyDDPZkL3El12w0uvztdAixXHa4xicw9Pq2Tq
Oj/Vctxlte3jztWNFZ9bVWEa1dEbKJK81VkBslxEIRZsaYfCC3QN24eGQjIvkSJJm4/wcFrMRMie
wSJzKTZNdu4JjP7ANi6QffTFh0MYHa+B51dxSvxthiyfAlUwrdw3Y0uUfqd7PHHr8RHa18T8QScf
3LGFEYgu41Pek+TF3T9SNaq66WgoX3rm9zr5hBtIx6gtqT9VHQ3SqGiCW5D6PVNBasZMtKDdJML2
Ehyk0XBXiCGIP7ikX+hrAh5mJnwD++yvMhV1pQuLtaGw2J3w6rIftYLAd6eXv6vZu6ZQtcEpSO9x
LzbCOV50xol7w4arTe4rHymfcuxHwKsSVCVzD7JKGzg/LIciTJ/iGf1eTZWpPPLXzjwIRfdVBUIr
cARCreybp4paJC1A+ARpiuIox6HtaPTzy13ygdkOwSWW6Tz6w2P/TfGq1ZzYwjiX/CVmqfAC9n/p
kLiMu8pOKYA7cCVYgEsMHsOIrlf3t+bmUE4v2Y7PZjbVDVvuuUgOYffPEmgyfYchHBsp+oEE6GJB
AN/6H+5k7Wv5mrxRSmopjChm+c+XoIUq/6zuvkrRQNEKk2pcSw6f9L2shk9rwTbrYLAp8zx0n2Do
Cs7Icxyd1PBv6NhtOkDeG9NG284z/Hi5mpVFNkJuUtLT2+A833C+nrN+Q39MAcwmJNT9C3OHZxiH
mtnwsS5fQfB8PtsmEkNXT5VlnMqSoiR8FcGzb7/ejgXQ4vwDZv7fHOCr5newTC3eI778lmFF0JK1
uZvyqrAlDpGY0IHX5K6Mkr+lu96yp/3Z18MDEa271+raZ5WTum6TCdFCjq2H/nJ8wLc0X4B2X5W4
hWRosSb7/gQFZUPjxlt4T+Q7sWaYRsPqDd0jRTr8x3/jlwhEb+kNE2aPshDGSXjyjC2E0izP/JNb
H58+19nFBQCdsjtgCC7YEOI65ySG0lEqTFnKzrh6FjAzoYbanur/buOWu6Q/1GScylTyNHIurnif
Cg3JzeHiwru1JBAoDeogir2Jd4tYD60lXMqZci+M+WDLdx9KEB/o6bDiqCb9uZJQ/VrXT8PRkBRC
VugVxU85PFPPuYBOI6h3eefTadMeNsKINMZPpLu73IJtrgJE3vCh6h41uTdDZI1dErGQjLFqXTBi
Et98mFnRk3tHHmwThlRbB1+X9etNqBWQI/3qm1jSlTVekEu/HWKwosrmq3OnySMJ/QPsiaNHsvWX
MZx4Ffo0eTJnGSVYpnys9IeQ2hoc/KvGqgDlvk60YXHHqBdbVS6XPI3p0jYR5UJgvlQJrBpaTG4w
HXMPXOCzcXp1VgoJ4L2VpWc1kEYBGSaqegO5jPmmZi2g+ENsIlzK0GyFJOetEoEgivWXGlTQZb/0
eSLc0yMJpxL1Hogj3I2SOwdY1dMw9OSdi9+x3QagAZBuKO+AjW8TVA+E1O7WiwmggtFHRu0lTPAo
1hgcjAECkqyMdRAhG+zWTf79Hx3eDew/Ec7c7JDVuor9ndoQNrEKHODp9UchtgJvsS2ta9zIGL9+
TJuZcJSobzr6P5gWegcKsI3GiuGPYd0OGCtjbqpJqIzqmoWZJXrzBtylQHBlBcPb64rce/Z58efg
ulyZp1MBz7imPWgm3SkaLdAkWY7+E3ZqMfGQesVOkzfoNNLaLGDQDN/K34LHO/cWtg+EI7QkWvJe
wxQni8AZ8eyN9HHLT1jJzBac2VPGZ8zkGE/PrHezgj5Mic8WF5nrHHF+G7TnxbV99qAJInUkkPQF
0Abqw5M3ptr6NTFm0BSLoLOPwZFpU1SoOuVHzaCe6s/9KdctW/1Ikk8harzkKsw6DowHBUFenwkN
gpaFb6nA8rcATxkFW6/wFRXs4yCNejjV5y3qW9gNpWiBxlGckAwNE/lqF79gHsprA6zC8cqRE7Qh
xd5eP5P1k0q5gkdorGvoRQkMTdC97+iYldTzWKU1n+kCDS4bQBlFUse9ZF1OZcvsOS7Ixd7xbOp7
bvLb5rRSkJvoSEV+MEKW93vlL3fipRZ2Ulp4sSMF9wjmYXOpGt4B/XE/yZeSEWL1iDRFjyFEdrOM
Pb093AbLopDn/tPEUPnvz++iQYt5IWwEu3MoA5PnXINZ2MWu9wxucamQ1Y8xORPOaCy6TbIm5pjD
WYjHROntmaG6vN45dOyXx+Qc/jD2vlNxIwd22FJe0YYKoqeO/JnWCu6/n6CgfZOolYTb8U85MvQL
HhtYeub7R+YLkPjP2UZDrljvZcvQzOlkhuK2dbUQouBu/3zjXXvRulTct0Ngc5Gdsbc8deSP8bSu
TDiu8X0ZLX4ExY/8yQO30/UxM+hStF3ZlahsSPHbsv2FOY2/gDItu9ElX0CpiVmPDFF+Cn1ZtWOv
gM1fo/LeKOjAWmA0iDGyB7+SG3QNJi2FLfIGFWedQGv+duKyd5yz0Ju0dMimyDFxN1Q04TS2PkMi
9BZRpgtOXtPjFG17LPe+eAY/xGHaBYUUC+7kvjC/7coozGdgtDgJlWva4EFCBJWpRrgmNbofayzR
CRvqAVz1lQvtMYv42eZtJFG5ntTM146RcbVaE1H8xOlGt4gjqpH59mobOw4zwsE/YhyQbAHFmpC0
qmRkxBpepG3/hXQmRnVYMrBcReLf/b+QAr6RDA2y31BUtLmuv3JyDdBYE4qD1UIXcqw2SievQyao
st6ZqkzNQsKuVWQdzHv4D4qfMpE2dQjPTzhWmPrWROOMoMESDQfTcigCVa674a8J0zjE5yYHVvgA
CfTouatE/Rm19VgxC85Xk3qoQ+L15i9CTzOM3ykB4LExZPnYl+U1waMYl4DlVg9O/bwqvmuuam7v
sYpQQGv4RgHlWzFNcJc3M4nJFGC2G48ETNbSWqy7Mo9UxQ5qpM9LbTFZHGs9TJQFpg7agGulozMl
fiawlWptrzEZUgFkbygYoQvXV5Mioa5fSH8cNS5PhzEThmbjHwuan0fOVgE/bFgPQPaZk2sXOKOF
gdKOcuNQAKSuQQQpVu0zqiPJ3XqFp4BdxB3t4q6XTbM3soknxxwUaOS4Xy8rr9RxCnn0hYnY6fBY
R8Ybj6YmTRFoTHcKVuL4UgJ8LpX+dRn5DjP+WTTWVDMD6hScCQncr/CHjcuPxhouQlVbi0GBEs1F
BATpr5AOmBf1eYdU8TrJjGwtYRHmOtssKyBO0TeKUXavWXnQBNAzbOYH290i61gHLnDOh8Mq7uMB
Ho5VlHe6Njti0nwKUJSFAPwZZDQlEnxbYOqo9LJniI4Pm9Hk+OcJ5bfN2hORXnYOIzjNIf8ZJZ7Z
OpVw9aOOCVOxXNahynw3WCZl35HB2HTqRaj3zVnIls40/Hi+F6sqxjjrP/D2Aj7FGNAzdXd4Tptz
gZ+VTJt3Omqd7oZwD3NF7B44Da/9VkAQ4lq8yLIUsrce50jbDyw/YWc8liiaQ4wcmwZUd12VSxx7
UFpPYMuNkkkgeeOh49IgysMetGPRrnWGRqKS6alAYJSpWX2B+lVMo5Rd1iV7iPIxA9D4YDFD6apB
wQ3e8MtYCIxtqWKUOQy0OiK6h9PmrZ7h4RlMDg9m3VedInQN6tznJEq9kZwnwrMFaLmS//iWsK/l
PrfQ1EP2ONkS/zzCS7F+Hay7NLnCWm0qfOBFSNKCei6hOhgDbVpY65hF+WATCcQzGE3tV0Xok5VT
knRuz5IoqwcNX1FIqMI4cE63IOqzdFxej/d4gdS6n8jXZDcWTiHxlnWfLXsolmPbpPgoyPaeuItM
WUivFImGdWFyIhmdF5px8TKAP47v6n5LaBQ0Ed7kVYUM1lPR3COD1cvX5SrN8XJPK4XROWY6KCmp
RZl+1o8ekhixdqtB6Bv3A2ZYhQOiCsMLxJ1SjjsLz0sXuyMlzW/YrTXOey/Al4l/m5SxZTg4c50T
uxNwosjjAKdX3LtZWerNm/RBiLligZgPlPy+2yBumFmiCSvWmXijWZbFC6droo/lc5guPtysL5Iv
uWvXRvJL273PVea/xKrIawn1byZRNz0XVaguB2PwgekdUIWWiL1v+I4TMyGD/eDdKNuOlN2pD/4z
5W4gLTkTfaoYy/IUG23t7Uimvwu6Buw+C6XzvUyRgCo+pd0qxiKYIKKcoQJ/c33ae0ynIj0dcAY4
6N2v0f13HIUh6xR+Wl7ufC1Usd4HZQS1fSiHwt/p4Ie+G3YsW82cKnRkGMUCXqHs5LSCHvZi6Ohi
SGOQk72KWT8DlZ24IOy7Q2pTAwOMhxUVYyJhBDAhJgGGBDRONbqRtYR6HwPSmRdn7YKB41JkLcIu
oWeynTtnEbNtR/ay4oa/4ZJVUSGOHsSm73BBYYrDUObsmK5mAHmTPft5bAi2gVsuKJ1S0SC/+zqS
2HrI8TmMRgHj7FZhFYF6CjbmABejgQYVrblK2bbKZ4bYJxIqaGhYuVL5orVmUWrGWyw/F73/0C/y
C1zZh4+7jqD7k+UASHZlR0VKqjhMc6Nilj7tzP/Rm+5G4+e5+4bhFTLPxYjfRx8JnAH5Jfl1kkdR
QDNnRW9+pjlviPXH48hkAG52NVY30wIAlCAxKH3+W8ynDCKwea7I+HBPvaqrs+s1glJW3Awlfath
jsyeVwi7sRfRwrkZPnXd+bk5PNqIl0BcfXccaGSi9joz1tIMf/Vl4OKGHHZou7kmcstgFm90k1pZ
6B866E9vCmZuFAjIKm9v9/VwV3x0ZBk7mp8i7/K/bYPkYKDVU0Q90vngLcxs7dwQsh8O069XL5bQ
mwmWO2I3q5gAHpH1VEQUFk65lUiGTS08t0WWH6aw7ZnU75fDD4LGC7N/AEeuMFRg8WO7jEpUljUX
e5wA15HAcCN8/NDfJQeDkob4BTRgEGY7NlMv3MwHI8khqs5yWlNNtTVl3A4syOKxzNr3EbDl2N5c
/zeqQchIsWmskg7HCaf4XjhYsWDpOdQe/L/RGpFeQz7Fx2aPD67WIDtj9+UTc1yWjR+1GmaBW0MD
QpIvzc0c6O8TNMpg60sb/cicMdcaDLCn66f/+zqX3JoYUPXpl+ACNKfecz+k2jRf0ylc/SnT1SGb
MfghbLg/MR2jmCD1ZQDZm/WBr1bOPg+j31WhbgsoNilsgES8YjqGn5d9kuB8vQjQKV9Y/HpMUmU0
tkOGbMMIQrOCIOByGJnkGJS48yREAh0a669A8EJlX30w/8B3YHgRiWLlETvPgADAp9e74MnVskrE
itsPKCexAwW6s6xXL/4F7btxlShYkwFEetiP0JrwCVQhTb6BOSsLDW9DKJK48p/O34dmiyOVirjQ
5UI9uba5CE2D3mYoRDLrui6aY6OZTVXKGYI02I+6/JTTp5Yx+TnW4eXGXWtlaT9CSKqJB+2sbWlH
Eiq9eDmIfGpmc8/+3OhOYJsXOqaPKowEEbI2C/fnRnEO17SKE3UpRUfVhKOrPQA5W9UK/dU7J9XF
haBNfmc6rEKslokmojCYFxXRtrsErzPnZhKxOa4vBMMcQfwccJnHOu6lPhb5htTqLhLQxEgq2BTj
4UWqxN1mMQu/NBHNvsTHEk+J+MR2Xc6BsyFYe8E4ouDTNOqvTXkokTpTgN5Up1XrMS/Qw/79zxmz
BLYqUNPONm4bywSxkwYdXpVnzVTLvJLLmZMZ5Cwc8RCg4B1STHnXsaL79vS6MXd2AFjAZjuBpH+V
ey1nELM/z6wrLVMGRsW81Hb6VVxyI6jsz99alMuHQrlyPXvsFj45efVfSmm0GH48XP0KNyoG6g0o
AegAqGo4iAI/AuArQqgPLLQaLZcUF86AF82HoOh7JcEnihPLLB3NdTqLTvp7M1KE0SE0TBzoJT5N
ycum3/NOdQZh+SxcTW8g9pv9TQnIokkCQYl18AlwMQm6cLOloWUvcxebQtksHbW3lnoONTwusUEq
qS2ly66HZm7R2HwWzrW0arRo2VV/pbDX/GvhLOvPPqIzRqqlMhWJXGL/4qAfU47tUqUAesRL1R3S
W7RYlpuaPjQHGP9J4eXdYn/EWDvM9YCNOJIwUL6TuYD+ABPy+aJXSWuMoX3vJcb5pgCyCcJmstez
gxj0gXwGjkCPUNMHZYUpW1obt2POE8WCSBhrJbaL73N+jSnon+89GFnptkCRD3ZpyY0KaYjavHFJ
6eisQ7goswIUDP4mIZViFm3I6otgfGR7k+SbaaAnrFbAkv2l8tF7TLhSXJw7pNRIvXvuIvc99k07
tPsEvxpY2eTtftyCN69jZl913cU8BGpccSoEN52+Eso+WaX7xSDDg5ryKET9UHyVaT4I36Y2zJva
pDdILcDSeTIlinFA2RE38/9LfChta6io4rF0eRd+oOyOtIWMxsvErZUjklUzjULkMwmebmyH7Igv
0NU/f/vHtKPBFNYOrkTd2FRmRT/22wb3moB8Tj7yrwljC1X0PvNxzOEsd9AfpgybvDvnxM0E7MXZ
CXAkV9ICCvGgSizpc+77JkaMOIf2kyEF4uSwIGHthKm3MqlubvFMIc4dkZGBsxObtjXyAfEKwbCJ
cD8OWf3Qbv+mA4plIV7VEV/lcd0yin+27KIdp/yfqN2b43OO8EbIrg/C/L7EWgW0TZFKNgL/PtHw
nVFuxoJ7dirlulF3+efhfNNmOzbUMqlb+qzQ5Bzp9zhY2bPd3e88+W2x3IHehAAk95vE8+hElvTr
R5SztRydZCte28l3ElTXC8vNkkDWRd3kTBDUb3UgrCwNuefiQhgNYnDSMqMl+cQnIBvwsN75D4Tp
WPEq3kB0VfVA4E8/gJoX/773I8qS+lrFlG2A2X5XMddoiBSZCtEl/S6XeJMf4L8ywSqAcRUls9vJ
LOCE3N9DRrjPvJhTQ538aclD2iQR78sz6nUPBktbqkPqdsFIUbWYjJLI94w3RcEVyKEwbztuAt0p
5MzCatXG53+5FiItEBchPJo9cuRSkKD8wtZQkXP6ExumHkQuMUmD/NEEUmiVgmty5bnDDtda4ybr
cbqz0uAYqFL6qoFME/llHXJS41fuMmUsum09UUNSr3qzTQSYKgpwT4PiJ6IqWoDB9tJJKzplQxD3
UkZnoOZCn4+31iKGcc/1/aNaDVb/D9KwfUk+ort97eHBhkiu9OtDpKvmLqPOsL3KH+oxtf6Fd2jI
Coo3Qst6tIKnSPeB4TgY3b+VeRJtPNFvxAYB2ccfz24C8WrIxyO2TLYs7S6n0NdIP04uRBafMwH6
H906ExRkUixMw/DpC/27LWk3O8G2vu8hKRk6BR6pp5LggtPqUtWP5eNJ/sbVXbyL1QvWnpzypWah
JeR/EozJQTwEtQN81A1F7bb/YNQrGhKxjKE2GTA7GlRZMCTEtYyFc6BmQR/Cy3ehl1vItQwQRUBM
rKk8whNLrTrElKeGFudNunOoJJNKtFYdzrlJlFAoTCxRgciWgp1ni2OtfqeiubCePK6n31opcTxP
Qct64+7hxys534cRiNUKYfsKCgcSXhR60JQnllix1uZgQJ6eTMV5z1yN/zbPbU67H1P1dG6hEvez
52KTtNDBHd0YTzEXUz4mY7kXya7Es/+P2BxpWwfHbLeW+B4O9LN+DQuyubsuPo7ovb2OPuMp7JEY
wRX0XZ9p9yPYOMZ+260ufq1TcEiQ0JMvBjO3eTFhbkl6HUSheDZ1dEWeImcgIyL1w8vtl4q2NOk8
xtWt36ZRml96SfuZStaps6HqLHwcSNalVb/xVnAQTBxywgsWxodQ+mqsx2hlwSewkO/uT3bjXm3X
9Nbyy60Nv2OeVyVaxmoYJoqbm3P//oomj9Vqz9qCHFyDHO/ropikHVlPrNrk75xUc79AXN1rN5Fb
yPRnIDDpHLmnVNjDWd/kFuH3zD4+AqV5tKujToy5yFLVkjZVODwuv+ZgepbluICQWbOZlg/umy1g
SDMI2CSx6+I6/WSQ8RllZYHcUlCRYz4XGb0A2Q8lmSda/QRgfto6rUxDzYO4UlHv/RTTkPo9WpNW
GM4ToSaFHbN4zI0wm6Pj2Dkxcp/398s5FQ5TqW05Pkg+KzxIIx4+9uLKOV+7JdxddWx7j18qV83w
4UGQPJ4e25ng5rVVkoWwRHt6PHvK2p6Medv/7Wcz3w4ZmAOVOeJuybDf8Go3nBr+qosartS9CZOI
HVqzn/Y7P3RVlVo3f+vYT+UGW21tXkk1RI2ebcekZS+HleQhwuAln35Kj3pSbsXrfpJ01Ftws93h
IrFrTTjw0K5ruQdCVynvVJeZh/4gxkyBUS3kJikbyDGJaGp48LxEP0Su9qJ3mEQzktHNMoNXvKc1
vNuYN+ak8qDssaRkC4ioN0yk2XMAQD/zBVX4t8Kj+2eOQJNVGe5yl6bKOoxTHqPYpNNTJzp3LvFA
HJ7KOnz0cgZbb3aNnMPcDx+rmL/HCDKNWp1LvOLxmGm5Dg0FEa58g+kiXPAwIxElX4Z0sFTVcLjo
BLkvCq+H3MejXyhb8gjuJORoI8FvUm+69cO6aIY3bJRReLis0jK/be9K/sSMAN0iND7+cR5PY9H7
dHZVt19oEqz8monxEyjyzZgNYO0kSnEgVLloLTrMxvQh9bMciPW5gCi5uiiThuxdNZvNRfsAFFGc
FghX+WIV/LFBR+k4M/Z/3xsoG1Nt9Qm+8DNvYNx36Esc+LIPkY76VJdlxxoi64IPlhb29PTO1Upv
BtB/nq8ExzaQJaDe+S+sHgl0o8LR6s666aiNaSpX9MDHnp19fth9pSiW29QrWQnh7jkt9vRENSzc
BTw6/UXWMNxBgeBGIfJpv472p8UryZwwj52ukhqsHnoJqqTnQpEWdSrmhwYhlv5vS/lrDKEhF8gl
dLoe0HM/5gbz0ewvlTqFnM3oVheqxliIc9u7SMDYL6lbyJLLmbw4G9sZsaSky63u5vrJVxODBXVI
17C5ex3ruNInk3c9/X/9RbY+2GTdc1RPH2JgNudQVjbjNpLiHbZXntFR+WZX4I4HxoqIvtuf5qpg
gIuO2dHXERhu6dwv1i6JCqkdGrn7b/O3z9zgXC4uxmzi4qxYP8WQ4xkLh7vfWM8cMUICwmB+SS2P
+/qDK8e2muYcUBEYYCLPwExDg75n2FON0DJYdAG2RgwNwi9qOlL6uVz69wNroDmoM0Aw/sE3pGLC
PsZESaVgfu9bJnutdMWz1pvSh5DwGxJL+H3WJlWjcYVgMLnCQN0SFMNrsPjbUG1buIyWmgObYNWy
pEimHpLcB1eGQFm44pohU1IfSN3YWeoDzbtRNti+TUOE8ZtAb0VnsuRnzzZYDlyygB99ullBj5eQ
RcGu2c6VYl1XIKTgtw8EIt8gCj3GqBLUgEYjS3A/m8ejPhpUXz4phtFuTAmNP0bfsh7VTo5I1U6V
O0i3Us0lUOpAPtFZOowKeneeGYz6l0JHQMLm5/3xLZlKv037tngvKktrhdJ6WhAx0jhUQAhiKokZ
vTq3WdRJEuOOH/2Xd7QHwyIlWQW6gq3rpFeF/piYD+VNA6jR+e6HS5+vnEardi4c+/Uuho6ETE4P
tGnaHgxiEgcWjjv1M5z8J/dZBWTfPzSC9CCXvAQkxPPfa5xDhr5alyPhjQO+vr0Qph+ddKpboSg3
V2JOjOkhN71wavMUju/Kcwl9G9tacuoVF0uP8t1LV6TlF7kB6qE9gXDfrEd6nqkhPEbNIdPwSSj9
daDQOLqQ8D/juKbsLC1ZUBAiFYQh7XuSTk0DCwRWAj/mbTq6r/HWeKVGu1a5AjCdHWxjkmAWhZYV
sq62lEoYZFKUGYxTmtcn40UEMirzjSNbc0vx9Mrsb1yj0cgcOod5C7FuQMYm9G6DsHwQNfYfWEzi
iquiuILRCOs03UR9VZ8Vx0aUXbOetAWPNetsm/FkAFPRErunNhmz4OHBX+bm4pTp89glwMZUNAjC
yFQNiXwxg7CoxrbupF7jklXHezgwVm62Ki7GpEeOTmXinJwINZPIYIAGw8vGmQPqK5kAnVg0EkqH
CWjVvvLWsiZ0jZLn4AD/35IqlN83XgU0OuWgs2IZK4hbd2CJv6T+m77zFoKTcBDc5m1wI8HHyKm7
NyUGF8SZpOESHQX3eXJRGpi+d81lKAiio39WGXZMs4Dig8r2Kyim0oWTiqLe4oQ7hrXlVG9Wd9/x
buk3q5i6v9ro2jDZ/KJPXuDZI3bsc7jn5HHwb10k0o5iGXTnZR4CkgoYpfjBU1C7olKQq433cO8U
gBxcNiXSzB5YyUivzZmvFPqwTEeW0j4r5T03Z3yPjB4POBBeTUDwkRguoV0nz5pPyIKdQFcbCW1B
+AUpkJKyaCD1yvF7047S9gQV9oqlWyyUvV9FQbkmCsdGA0r/dD+obUGr/8B9XTB7KWfrRBhM/2m0
Pp+kZ2BfxpOpqZ53UrPFd8UMRSNCUzh/qOX3HRzfntisD/MqALC9hymrwszZsilIvMtY0xc8Lqfs
ScvCmwTrUiSlzTLJFcRPoBjm/BsQma+Qr2FKLjMxYf+EEPERgJaPXHYSiQdKS93D60zarCkyVhAn
UCJbbzxj3cRuwHZonY5E4ICOvU/rEaJXOulrC1VV7zHPfZW4Ewk+Q236+lkxSP0Sl+bbW7Q60dG0
VFmN2RyrICyVEoheNEdgFyqXpwRQILgIDCylVpeeNxM8yj0m2ogAqGrITME25kFXzGibp+jvI3NH
9Co1NsLYtsdN/izYzwC/Nzbiu+b9rrWMW/Wsa5ER84bmPFtDVYiRB/ar52C4luTDCsdhxZc5HId7
lsU8N5X/nR/ZKXw0bJdemYW8OZVk2PHOR4fRRQTKYwm82+sscE5WGhXC611fsEIGG2brI+NkDRxu
HpYWDceUP+KQNEXkxJB8Az1Mh2+AW5ZAk2BeBy0vcFb4ZmovtoFCG6QuZBa0DTs4x00/04jX3rM6
7cPUvF0c2eWabeleEt1kITVe+RSnjTcoNWAwZ6vi4vr5vW4DPMQN3okojJDh1lQPdySGu2Xumr0u
iDCtyZXawRck5P4+UJPLZv/go0M/Kca+d7WvzU28PUfeRdQTpvlg2sLHg+kk82E78gL4gH2v3gBB
rN18UdBTKRDcwLA2MTW0H+sSUn6pFLWsSGDs14mZPkdjrtdBOKAYgco0yG934IDmf6ZHJqoPxmr9
RywKagVZYnAP2kOLCBuDQ7uZz8qYqa8bb+z4YzTM+Fq3pDs8uDRiM0Vpo15K/qe6ZPxBkL+vKm73
bUTXTcz/+FHm5+UbRD7XAvr7jMjzI+DrMRizvsATOF42BeppTnBen9K4XQc3rFn2Q9FL/igj9G0K
Q7gs8yXge9MZYR5h1gM6F6+B5kihLoWT52E+JJ0V6gWR/6Sn3A+m/VyM2KLMZ3KFwybm7FwQyrVj
u+Dv0vodpYnGRQXE9az2Z0dAfp6w2JkZ7tdPH4wIY74PPdcXCBUne1abdjaTc+a75dcMY5JEbHeX
NjEdtA89sVOQRtGyylBAoxyTKG1+odbhBfaOTiZH7vidoFe7tmo4L7j/bA44A9gQJZ6eZ4TtFmv/
cwliVBVA4Mh2dhs0GgkYbEwu8iSdnibuHDxyfowXb/6f8Gqh2tNwrRujEVUPLzyhN1Ma5+QgVFlP
xDyHESHUH1SaHNxys7Z6Pki7YOAnhugpKhba3Vj6uUPqol4BcNDhpwnZmuLUnksHmgoQshNtRS+t
fKsWiRzH7AMvm+sBwqTas96UOKXf11UVcMz1Sk4aUnGCW+TTILrw6j41fHZycH4ig/i5YS2KR5Jq
ta+CCagF7Pw69ZrKeAq8DbwWKkjb82SjzVJiYSVfRmP7J3IClm00OuSQfF0QiFY/jGLjrI8D0eR1
kl9f2mson0XoCF6vAatSV2/Gn2lseImfQrUubSucjXBoEZj+8zy4ISRIgGwJIS7j/GrXihY+K1WI
WwLcOxAbcXL+yv1UhHBrbASTqO25l0yDqm4l5CE6QRpSaZFdyQlC+cTqYgPmyO6S6JhHOA0cHZrP
XojU0R8nvAMN76wbPrQCW497Bu7nJjBzv8evmbCg9A2cLlQ+ypiH21oX+lVTFfJwE479CIAImWdf
EEmq/ZhO6a0z+b1icvdt78loAyhdpylcRVpBQriVLehd4Mm2g/SvpCurPYuIHAqILJjdt3Njvris
z7JwX9rllB8b1neLIVOVap7k1/PqDA2MidZTIFfaY/SgkLTbs0WqOHieF6DR+06enXGmhUBTV+tO
2Iyx8VPUM9o6H/N5xS3z33Ot2hhCpmM4gLsCA+CmaVFkBYWVI0RPCZjuP9nARKKa7K5sqjH9c5gM
LfOIz1pcVLcHgolsNyK4RTUceTb1uqEFExtG9jalDmIC02d+4FaXzCko2oSTv9c3uEgBrU/TC/ja
eWEuqlJMcVIZZ+32tBGKQpaau3XW2Nk+H4yy7tem1vXHC7LtTG76j4VRRdg4W2RF0dvKdYiFC912
h/9V/WkphFwoXFZKn4W8ijuXkOWXWqgLiE7W/KmD1we7zSD+3CtFR/WOl4ws6nyBa6ov3d8IzcmP
yrhQqvZIM0fJ4qvd1ti+/qjFoJn6ps8J3E8Cpxs2wCiOX6dCDpHKjnHm0QjupaFotNoI04ROVaHV
kU011cT03GL4uhCn5HO6ng0XSSfLKuA8jQAeWiY16tRJ4xwhCYx9ch281fN2ZNoNkyPYqNmjX6eI
M5GVc8cuZvhAJAYx2j1FPvK/5drs8X7ie7eLe2LltF/8k3RbH6OGQ31vueiiXZTCBiIN3mU5nUud
H5ccsNwEg7EHZy0JGy/e8TRLQMB3K5EYXZ+T9rt/qrdBcIYR6ZLqlHikuJAL3HTs288o3urr1pH2
U1/o/nmz/RUrO3OwlRKaumi2Tz1RnzIDz4Fed3d92/7U2qQaXtL1eiulrg2tDxUKRiDZJfBHOVe5
SH9pgy1HFXG1JZmLTS9Yp6GfieUCoHsPhH4MmBpCwMRaa+UuXd6+nW7ZPb74SQaoEoJ6FcsvYQF0
SkUnpThlVRKGrK+zm190ZWNGBnbtzEiTpV6bPcu3yHJMmFzEsgzfFxd58uO7m0p+rXHMMCMzC4To
07fRu00dXuZYlV6L8BJUtiWFta+Lr+5v+lRNdyEo9hRZO9R5k66gGES8qNu7hmJhpnwA3s3+Tukh
kFSGRuVTecrTnPVhiph6VmxIQLR7IVA4wRTnY+5ce2unNDto8Br1Q6wfGZBo6FosiO5Cfe+xyKnX
1DyTmlifVNXuuRipiKhLq7c3PGgSi51z8Z78bgTg9CoajdmReJzxPGTuA5NOwLLw4+/6Rw8PkDYr
O33IjSMJjvLQPDyOQ0Qi8BWn38lcdR61BdDRmSXotmOHgtmYgRD/Pz1/qi07LKjIUwDp2orl3maM
rtOpX7lcqvDVBzdSGoWtRZt/HyOJBA2TV2vCpDTwMTNUPXXYofrlxsF49oqZt36mnwSNFRIW1Pnm
XiFlhftoggYDjo/RPDN7eqGevWAPWbcXYa8zvKD1AtTTBom7slHE02EopvExeDPnAET90+8Gdxh4
khcEYPhHqaIolbT+9WDkQ4J6469T/Op/WPNUh4HZcH7mXaqnIKukkdd7nN3s3XbT4KJJATVf+u0p
xRil4JI4A5TB+RZ95WVCP2rQaXhNbymKsyhD6LOKYjQYyVgaKG0UA1T3CGCc5b7yfPn2KBQDjjnG
aDPmdllCCXIqADfZp3cyF+uh75FdOJGUV3H2r+bTIQcoyiYAet0fAkF9Fy2MRN6cy8y6aeOycDnA
/DGzq4r/d9M0xfnavaCwa1biMfLqIThvlR6J8OAczU/iWtDkqpUgi2LVK7UCTU0AMJPlV8EIOrcd
R7NL0xrBxKcdiFdb25rknO3NkN1uZgFt6Pw3dFHugioAmUHNY0s+/qtUG1Ls0NJOOl/xT+6ZTDzJ
0gSU6FJTYpMtIsnjUiWbiwbfbn6f6z1wCEdslqAxx3mZcYwCL6SalzsTiQKr012u8tBW+yMHGkv4
ZNPxNkjccIswHciRghAsZHNP1FptpUb3AoVDCbNrbQbux5NIzQRIdUaDIjPdjd3RYEtQcvgwwCFa
LpdxsfU4cUxHrZqQjMf3Qlp938jOiBTExgxj/E9ShDYaSI+CKCefX3apKl1sA2WPMIuQjLFC92Y5
lShdQlx2Q+FkjPE54Jv2h9miKCjGrCkcZFNjvZbqwHV9kP3FJX5UwlD8ltfyop9O1LgLkqWT5qv6
wpbV18I30Pv0jbKACQP6rSNeuhw/b9ikv6QUlNXOJsotmrlfM1D1XVaBou1LI/sRxkUpMFs4KeXz
w+5NgkTSgqNpGwOVBq+HrI7FCrammCTddmRL8/Pu+T1UwNpvdi8y7GHnqIg3zxU25MlCY2yZz2qd
RZI3EF0v8Fw2v5zbuP6tVeK0hUn5n5iDzat+6PKnxiKXzTmu/9/sgWREnBALusTO130ezlas3Rp2
PNqzvde46d+it5uvjtsNLPkHSt5zrsI0FSvdmqrKfg0QFglVHiib41lCvN4DGb488DtZq5jnlPPJ
BpVnHnKcdojHIGvSi9FEtRi5dUL+NIH7vBCX8sADYgOvmJjCFyx3WPJMsmD2m5e91l5+J3kIK/ii
FtpF0zheLRh2rWUWEv33A4a4Evm3U4CIIA0ZC0vQ0bdVu0YuKic4jxQDuFR0VWE4yZuFUYvpGMhX
fu77yMgjr2/Wf/JeJxKYLQRE9uACs/PS90if5CLbKpFOgyU5A3GGr2AupG+YGcHiGdTA3sapI9h9
zSbLMAftv3saJIeXlP0inbp6Ux2J/soW/RgAc59UmNwJWU8sTFBSsg7qvPIbK+6lcJ8TvFfbQFGA
75tuubTH5bQzkDcpRGB0zjL86rNNxW+3XdJpWf++/rvJXT9LJj9T25Inxh1ufq0Rd+J8/gdo81W/
pNc6ONDZz2fznz8Tgcn1IUwETeIjEYfbOws5+acRaZdMtZMMjxpuUWveMemSpqaLXNruKuYS6P80
LNj8AERm7LgRIS9beTsG8eg8dZT8wANTFkEqNaMyAaSgkf6vw1AnO5dR1aLjmHNOnO6RRgHOGzuI
IHaf9JN02m+sZciLg3JiEaB/DcX30qDKH/O2U6kW8e2bGls45t1P5BUWW4Rlsej2uHoyw2Kjz3B1
hutdtxqPLd+Wel+pth7CobqJco1vYNWyRxbilHL74oDEeTJI9oWYCDfBwn9yxDzf9BHsxSBr0jtY
7iE4ci4O+S0cbW5f8o4w7NjvAZPGzM0n9W6392wz0SqTvf41O8iSQpeX0ybVl64tDWoK1K4Vze+T
0UTv3hgX8gZiICBbiQTAYhTgenqGtjDyD4c5FYy2km5rC49NpNCh8qHV4YMP/zGi9vSSVjM/Hok/
CdxuDLgP3JCJiFvcjew90JdnEN+yMkUwxZnFl/VFgom2dDk1WlFyCcWlS1R+mh2sWsTbwdMWIxTH
5gBc3/IOJ+61MuGywkfokkoAQxoZ+Sz+bqKFOodj0mHIfLavkaq0b/ABskzJ4+xNZpsRqq3GVs/4
AhhBEnbCcOXZs/BbZ/hZBUU6rfBQoIib22TxOQaTdNxyUml6qXnoYPLHfoY8eEkUyddeu7a+KMI0
91OhNrUL17yHrrY9MIaAwFDOZdqJlC0ZoI4y1vdZ5n3S3DV8/SLbBHBQIuhCpg0PHvtR1eY5x4sV
dt5eJydkJ/eUzzTEtPu2L+h1C70GdcAKwOUVH6AzMKiHro/bhQB2RvHRdCN/gRVFnxqZyrDYoYxx
lwvZ4SMxFBfe/SKneaj5jYWiF0iavum/ApGgLI8GF/YZ2vwI7tmcUk3o48v1l8NJFYY7y8jrgbz2
KV38wM7VpSpDLuvlXslRnl9qptQbxyRaALtF7GHcbequVDRVf/z64DcX+MpZbHAFoVZF3PbZ9AB1
hLnX0RcoLaicBOec/r5gNE9UrBP0Io168F8dcjiBNCbWjuRj3cneIIyiSEm3EYw4xMu49gbsv6DU
Ydoim5ha+DX5lT4w08jLC8GEwML6SE0pqGMj9PRKJHbDnTW6u7IwDvDiT3l8jsJTzj0krbJD3xbB
0GfAWcKhjoODJVipCpyx2xlP/o97mQaMJt9puvqtv817n4zROUfs9q0TBAWim4OC2HhIRuXT6uDO
qMaU1wojmLZMXf7+1jYMuZ3g+ovDnFWwT/BMibcaxd8btdY9+/pgBmaMgnZuEhMG5KmwzUbKHhZi
9TPb6E55LyyblEnRyjumQah1Xa3vmsRilX9wSFidqAQAVxBrV0HsOv0ldTQ2ZXZ7KnvcKCa9D40X
XJUyVIu2PAUPzIg5r7zWBK7ILuqFnj5XwJnoSurNQohcsJWHJ9OnEo4lkTg2C1h2IUFdevadCF9t
VOtfh62TrhaUCeuhVODkMzf8qPG2IChjrAAc05C11pd4OxvMNUBZ4fKKGsJkD/iFP+siwPqh2cMO
+VkbNmH/8DMF8JNS0KlsHLZbnxlHJiVsApXCIiQ9txIGkSVIrjbMqbFed+yRBTvcKeJSFLMTtGX5
5D2emoE9VB1Q40uGFdpl/Oqh5QauyFbq30SbktPZJg/xjeuqCY/d+SwmTokzXcqol1dPzKKX17gk
YIgC5d/MXyui/pLvvJLbF7vvQ37zo/sLhOVjNn/DkPNu5nT+Jhn5M/qHcZZy6yvRwZ0igfUmydm8
HY8Pjzi9QamZUyRRUy8BftiJxIdPJoeq9BMuIuT1pmBx25NYVgOaS6A3WdlT6cKbuLl2zWcmQKOR
n9mDyztwCB4AW9rkRRFqF0r8zEs38t35USTb90Bq5gPTUlWp0iVtaYEyP3952GP/rEKIkkez2yRP
v3u5mZ/+Z5PaY/15Ni7Okn5G1lkJVcvCegl45zbjrC53R2R9YDlseBR1yJ+5RHTy++nKhJYdTnkI
C+s4GcSwKaoQ8MRVglGmewGE98EuLRwNoVgkQAsGhCGvXnnfe41SaeuH+w2+eJYceem/ymDO5dte
T3rdNm4SVkOEfvVwg2QDZqLzPSVE048xEnPanf2zrOTC+keMNeiUPF6W0dztSw++zoD+8JtNh4vu
+42YfegaXEeteqoRYkMw2j3KCCZz60TV4UcxkAUH7auv8JhMixilr1KNAZbXhnHrJ1s24rMKYxj5
LA/yksHYsVhszl9BBqKsf2xRAavec/s0VEXH5nhKg7if+ik+l8P+ooGJrrI+MlmmHXHeOn7gVNsK
0xxKh4JbN0atzEZLvTkoe3Ljb9eL+18r3I12uqc5+HirAyMbNGKW+hUteObK906S+eL6vMvw4GKh
cGR/SQs7rQ7/P30AU/KRTawaeoI73WKfeTbV26eCZzssvI9wAkkoARDJ4DE1BE60l5RbkO7iPwNt
Al3lBeXedcBxgmX7wwqhye607RFLXKCoq/Z/GKsb4BzoY8570+tvugzAbXlTinq9llvdJ7AAKboM
NrPhn6BdizXcb7Rb0H7oQd6vQBsLIFMSwUGPZEpjuiQIobymEq8M0RETYaYuW42N6kDQv+e9mTqZ
agW4vct2n6OOxrC6SR2NJKCSBZlrtrSqWsjXGWS5+eEAaUIocPxADWEnzYX48uIj2v7zCjsGGO5h
ivROTQBg/X+WfU+q4Ub83NafwVCY1c2fuWF4MuaG5d6anca1hEFjFTCf8OjygkYPEN+XTFEqgbsr
Ex0kF85G1oxea5EY3fpvzvAW9wD3n80bQMIEOCHnz8BLL665bicAQfmahJ8GmeJ4m3PaYbUyCrcw
82Gl0D4RBdWiJ34jnmHThFPdqBJCyaYlRmSCpvPsjr3ktuD0CfvgQ6sF38zYiG4owgNxEzpfd1LQ
bCoW7Hi3U2gomtORm2XGjvP8fgNlIP+HhLfkZIJV3b8l1EyaPn4Bi79Az52qZI1r5XeszpOKrkBj
mytLL0hFFSCCh8n8iEKxF2dXL7W/f+RncQV8a/djtIguBNUF+9Y3ZFDwAdwoOND5MqmoXHoi/vbU
ks8+3TlXyX2x6rzcCBh6MjnJNjHSGvS8SbLUMCZzmXnQ70wr+oHMEUcdNeeswdOfSw9YD/TfTNLW
wZol2rFRVapAEWo3nnAFhHMg+L/5ukMHyNj+WRz+cv7lw656KhZjI+5d+Db8Mm8uOY+/wtd7X2wI
a4EW6gTs/S9/7FVi43okf56zu2yB3ZUTcx65z21V/ZfSiY6YB70zeCcfB/jNBrxuOdGYFDjPgqFZ
vrSZbrNolid29oirmVeV4BHCmjRgn37E86f8NZ+8b/5B9Bx/rkGrO3I6WgwV1f49Mcyp46v6ydTA
2u3+idhK11NswJoGEt6dYc4tD4NFd9IIemwjx8HgM9PfqSuLyR/8jW3E7etdj7uROImWWlShtyZO
YydE/hy8VJUgFzuc8+tXX5aa/ekgl/6tpDxX8dbZxJjuwKgPZoRQ+vGYO/St+9yBapTMDtCaBeTc
weSZyio0N2w+PaHCcrlhOgKGRXsaj7NIAegVPvJk1JfBtD+gbhI8QW2q9UfCM8ica9qp3G170VxT
n93NLwDyad35hNsxkc8VgQO/tnbl3X5AC02Y85biWR9DPeVc4guCn9a/rZfzjKbRXE8ICRMpWfCa
sch0c1md8T4BNsWAQ7Bl50pMhzqoXrQF2KsePYKPUqnGrEx+3d983GWgTj5HO2swpefrQeAP2hhH
6PM5XtG1kMHYUuPqPf2ifzFpHf/o3sEMSPIT7akyvA1+NMU+K06PO+x2MVhAfaEreUlv514XqrRz
xu3YPN+7rLWLgn2MdWhSOhbHi+gs54pwwvp6q2g0fFPq+18Q6PvAea4e18Ft7xycGYp9sjf/nEqt
GVvaTQQoqLNvGjzT0zcoFzdM3Cah/WaH9kq+KLP60DS7r+RUhwVq4cqfeTP636azkUl1SQaDPa1t
Djbbqy9BhTS/aXhm5xSRo485UgrcovtTeuG9fpFOQ5VfJoFd3u8l3sRL9jg6XAL54JR6fl/t4g8V
Yzjald69zoC9bPEbzyV7H8ScHEbKsRTB8vhsp3l9Jtw/NHs7LTfd/93Z7tZf8S7oX0CQboqdukED
iz7XC6AgzM6ZJ7GRMUwdphwfM5i73CNr9upHGuQdcgCaNJqX+WDnQ4N1mH3WfVkMKqQL0owmBvV+
tHdVP49eWS3WsJNnr/RG8DFZ/qSq+o41AwVPFgDMgtyfEmSRg+/k6rTBiMVXxrSt/DupTqsIWPED
inoHt4cpFe8leF9czLiwBwCbo1bQFJKXhDyu3z56u+tatIRU9Z2hB6rWTh+uw6Zn/Zf00KgfgFKe
o6BAbOXTwH9p+A5pBxI9a1yfFn8mXuPChw/EPEZgItgkZP2+Mxoh/fiRWmZgvi2b2bFF4S3kXYVa
YX26a7QiaM1WZd/Wh2HDuLj+MVH+dAgw+/RWmSTUCuucAdH24mRNAfb5wI8HeSUqpZeVm7aaHLQq
RrmxelHkQsQPBNkRDn/1LVkgFxUxNOK8w3alpI/IAAkSzv5vj+WeIK17eNTWBlCqvFbskcbVixrM
+i4wrTLmlEFhM/BWS0PNmv3mRXI+56zY52WmRvtlEeZrXJP1Xo19x12X9tfbPKbfb3skAY1fpmVv
l+tROgtgX1LkzSYvUk58+91YIEwyJ18QvcJozCeyQ8HtftaduirbOnDddzn2XoVWxy4QV4JnPE2k
HYYmd3iq2++v8B4eoRFHSs3OCWo85gPQLpy7qBGUazkucGInM14piwfR+ArHQvAtnBzFiJ3Reze8
jPwcDIUbI+cyJNANTBG6DyHzgSuQb/PUnSyMQaL7cPKknszDYUQ1eKMHgpMOAnZruSt+x2gD4+e2
rRvJJ9o6HzPf8jBQd8JyFMB/D2U6oEp0nJTbFTxFCs1DnOF0GMPapairbKxnPU61+UQ+w0FVi6S6
YsuIJwGgnb2l7v59hSeXnTIDOE9T8d1rqkURhVYZOW5ue1MhHVCHJQA8orNfaw+P1fvMMFGaXMvz
n/mymyJM0+gfLputA4dXmxelKzEqFx06LKc/K3l3Rt/eYllmmbbXa8xyHzFveK+hTDKqGm+ka/gI
RKYY17u9hV5Nmc/L6M7gYw/jkjqJS9a093NvkzDdP4rhagZPjyR9WtPgc0hz1gUBxLNoZ+D6VJIQ
39vMmXnHv8x/Yi/Pz65daU0rBj1ao7203PnoXfoKC9fRHgBQBK5TeT+7qE4tPG70G/Ib2JBNgIVz
C5dYrhLaQrdhb6l0v01FL8SLarROlInZSwxEpcrATM+WeDaEFieboAdlTKEl/nrxfrvxGPgsWzH7
az23VWf3zWix97WO/lecIo/gj599T00SwGnwyuOTALx5YzwXPrPNliAWHj2lZ0bJ0S2VA3ZWJRvY
vLVasjDcU2Sw98UMgomVQpG2NDDjsoc6NY7jdCy+ljq0NMmucbEe52TJD20MFb/bymR+V0rFQzHZ
Khu+X/uQmbNZuCD7qHURXfD/018+q56JzVTv5F3Bm9K8oZW9aJKy2BRUq4pXpmNfelajZKwLKVAj
TUD2x+YhhibCiQtLn/UPSAcPOFtu+wWH2XsUx9PDO2euarhPxWimA9VRF1+k3stjvOLFTKvQfUVL
U5DOueRqsu7qLan1I5sPib4+UBSJ59xrfsuQZenVUD2NcoolgdugKrVrYvcdwEHVNiZnrJpNu2YY
3/zMiHA63Kf24mXSiGZc9ea0WJkwY/TZSw5F5dPfsEqlN54DOJ6mpG2Hy5iBMkUeawU7Giy0o8rK
qz0ZkuCZjQHFmJeorETHTUgxEFfJ1pGwpxCHBE0kd+pQXGRvjlofdUX/T1ruH8yjOiQWYPQSDVuv
IhodyPapojNWHX/BBLcfvYbj0/W+FQK5YjDFCfYA812Yw9erAHzN3hWvl9VT9nhTNo2KLC6PauJA
G8E44MFhAwj539bv7eDEvtQVo/hCyvX2QVquNVGb9p+e82BUq2xPxGuPLtJMsx4qQ5J4dRmGvs0z
KV4JveZCJaMqIS/fLd9xNUYlgjZZp0CIH23isUtocqY3qpiOuPQs+lzOg36UTzT4OA5he3wI6clb
dKcPVqdrmf3WQHA0ZKFWfx4RXy6e0c21gNDs09e4/HvjsUmbs7HW7GL3Ejy0yHxFbjCF+NkDIErb
lLD3nD2BIJHVHFnJdcCFZA3/WsFvamKm/uZ9ERErD2qd0NnyBTsLlbHyVnNUYrftigo1CAq/4z8A
EGnbziedb66HOtaij1URfDiAORqPkvyodorVmeAZvVeHSjSl5Ff/WIguyBm7+sz1ZRNwiRQa/jns
KrbmRU8aurst36ANNNT7SC5Iza9g/0/BsofZT/6uu8z40hdR6KSePVYJ3qxEq66lhrNQmicSIPA8
HPRMOUizHHkJHxheP6J/hWCrqf6K1vOEf/2QOUYSgIwIaTX30uXDkbi/VMj4MdCzU1U5wHKt4j51
VlJmxzmoMq4bRm9UO5Rtm2Xo0YcfJD0MRlSKpOcda9vBdE0/u5YnO9C0l0xDL29Gj0sP4I4uZYJD
13WnyI7OoYYoi2q34ELmnA6/U9fJiVbvu/U4LxTx7suSBqK8zYAAWJdohTkb6KTtJbctSq048Qmy
wdiBYTJAFXyHRPGn6lQesHcE39jehR1FEIejCGQaupI2lJCF3RwSI0k7mtfN2KJdyV+tadHWYLBb
ci9HDqT8xVRNVpO5vv9ySG7cUXMgUAxNxvXk5z9ShPlxcA4fqxONq8jPPCO4eo+m+tEVkQ9j3yaS
QqlzK494wGlWdNI4alqGsnUxhVMx0F41vn7igia7azHLNcQy4tVI014WV0Yf2kJyS2aRPa1OQ2an
DgY5KDah++o7SMrbHIxwCbqDM3X6tI1W4/cyPP+6l3AhKWcelSAfTyfdW+2T8SNoBtp/V6zucmpZ
CivTBi51wCfgXCKbICFkc7CpOBHDsBCGqxGTLOtWeaHV8etrylmUxZhTqizu9TXnTeXFHaT9Oazw
jtxN5kKQOR58b3ZkzD9EOE3B7zY0YFF7RbEX07jZl+Eh0kz/xxl6ZPoHWiUiaHK3prwO29SBxUcI
cKkCeNsdIFCNF9aB3kJEboZo6rxN/cGw0srGlj966uAp4VYPUV1LmRL8/IC4Lvm5CaaN2RJiWOP0
/wKuf88fpQl3D81UE0iarTLilGZFDjrhNLoLSWaPHpBJ8LJnJ3VD+W0P8VPecE4cJ4rnP+t36ZQZ
1rXGaqi449VTJUXG6TxTx62XcRKvL1JExoW5kbTy3LzIuiIQi44nX5d7xwRYm8KJsbhmpLsj4FQM
G+DTb6Hm4NKzWbWGVKUGZc0oqIw43N+hwA5SPwFWBc4bmCaVO4cb+YB0WsG+8dUm6udcsA/YhQ1/
xtPDHjAVEQ/aScKKfDq8Dyj22R2Yxr+tzaPaPEcdAD4ZjkH0CY6znyKEdFgUvlhj/29f/Hoksi7S
1ZeJh9wOXVO6K96uCmavzj8Bqr6HJeOGa02rKWqUQUJMHRFEU0BQ8+Po+mBUObGT58G11NVnCFow
oTKxyD6le/+mn1t/L0yRJHFhZJeTu6qbireqgdq4HVIjY+2Ee1GkiCKRk7KXPLQxfUcZ4C+OM5BJ
deSih1/FovvGlcupYTyqlNrh3ZfnPhkJNqIllIDjtaulp1A6AlIZNG2Iff65WpvAKn6CFlyNS9zN
G5ZHkQt/HjNTTu4Gq3yJbR7HlPKAAQoNboQrDgpWg7qkQYVmlBtWBdcgW6EyB7t0Gh7lDUzePsN+
sqiHZg7BhvfVUEzOrwu1b1YnTMLL2gt1Ccd9Gmuk+sgH0nx7a/mAaQVltzfneN5YeePBAq4XV53Y
kHJCiGlT0/4R+tKWHb5XmI+hrXFQo2ucaR4M0zEQvDZxHYU23P6BQf9x9B3T4NG3JCOGznrhrXdk
NqGPUZ4LbVu3o+dw8cpiOAdqkSJ9o4tiBkdTRakQAxR6W94LQ52Kf2iSLMNMRtm+52I9nPcB46sQ
BaaDFqoV4zvwXOrMm0iZ4THT5bF6v2uafgFKkTp6nNjMWB8c8jpwYCIN0xVBweCTHGIuAYoEH2fT
+ye7b95ZIwWp+rgh5/uDYy8bXZXVzZSg0bvTE9RKK5ZXdqK//n4oYgefg8PwzXaZXGURmC6ZM5pC
r6gCkrfQk8FxuVULy8umP/qaog4/GZzxhC3s95cdt6TEi/UmbBAjwQG2NrYusLzJ+y/k1zuLowsG
onnnAq48md8qK+qt7U7IsqJgcFbGnw6Eo35RQmF0lV7KwHnUePQdLMBSGVz0uMgfpDk0Ik1RfgzV
RAPTNsFxzZ46cQDudMvzg9A6ExrUF29PVsPaBpMe3w2vuHq/q+HoyQMc6/SCGZeYO/9iOtZqz09I
VuDoLZ6CgU1zHiE/2opHmwpPgZmRNA5itJstLl1DN3NvW5Oa/DQrqtZYxv+HJ/+ljN1gaS7Ulbro
EFg67BhJF3HXYuZuXMK4ue7wb/orYdhaM3lZkDI3tNQLsNx/kDUDpRNubSg0wyYDRMA91Ruov6fz
j/MzCGyAYE4kkhS4N5v5rI7rkCxsEjc1PgOEgNkguejez8CFnLAFB+66KsmpG8sjITNPbcY0UqDA
5thrQ1jc8VgQPz9l6BMaoKeMlXfOsDjpSp4vzslxEachvL21Cm8hrvHemLy9o8pE3v8cN6uMF4qe
EkEONZbnJWsfcchckzSmsGfVKT+CPb9/qapKWAc+sTTM7YluJIMRvOUOg513vSaxAgf3cwWNKp9E
H91PJyYOx9xFEhwClpn6M4Hp5Kls0AyIJLKN8UFMDFegxf3lP2q1iHm+QRWaHlxMitUY29kypbdc
kMtEKphGCDHRlM7jqCpJYJX1MG9nwXPity6bNRoFVkMVPYQZj1C9ahEmuAzoOBA45nVcve9cyazc
05MXIKBclg+mgSdw1u/IFMZnPDl56p4zO44KUYkQNe+vLQfHrLYeZu4xWTuhWtUkh6nxfHlmGRdx
rWbBPOWrxx7ha19WNljW9/EDJa7Fpzn+YM+ilYSlpiYW7o8sw/btwZ/52Ww7ArImKNerld6UZK8Z
HyCcWnIG4maCSDljcbuM7V35eL/3rlkXgo6G0In/bmOumA/+/Hc7xoMLzFNskdcQaXq6abdYH6RZ
Qf/hA+EmVm+pvOFIp8En+1nfozL2UIvRTncpJ6ioVkRrWWy4JJSHlbuJA+moIK0OKtUuIGaZH/N8
4MiAvckBu9atA87qCtf0HlVL5pzj1QZxXsJfgqq7u/yKpnZP/Pup3dCRBeBh00s5lZKKvqB3cowx
B+t7VXYf3jUFW8Wv0JGezUJNHlLdBlZjfDnD533Iqy2JX5iatygLcut2drRn9FQGFdyCmAIjGpUT
byUCAh2I9ffb9PGEC/5kfwSSxN3AIBRZbpLKX9PnkBbtNOxGq5QSpanblennLX93/k6WqPZky9kO
XRDzjlRGDbHHW+YyLS/Y08bs8TitNx1tGcPI2qdoR6SBGJix2b719RNHb5hTbyjRCrjq3od0CGN9
LRmXI1t/J1mmAPrKSc/NfUG7FCrJXfm9mdvZDsIiZL0DpPMgG3qOM+bPsuyIBsT3Ra60kOTe7jXF
yx6fePEhCLPC9S8iR/roONoPwU3SqlImzibwrkXqgGlJd7sYxxCvVQQobGw8Zzue8hswTY11BVHN
jjU3a6Dw9nghyqZvrWeG5aefCcysx1IWd1m8two8IC4gM2FBvVZ0fw4uSw0lpBA9e8nRXPwy2SJp
0Dll0uoRhYvJ2sqG9hVQCA/FjlJZuCBhLwshSCrtnUNmBF3jLgyl3SmL+Gufm1Ke94Vn2rzZ7S4V
oEY5CHSurb3vRxBxo8OfSfhs3nekO37gKQF9/BK8KFY4fb8GaLGIHV1XFGNWMyuzYu0ywfrTpHi2
J8wZkoQelapKaZ5e0prXWNGIpA6AEUb/hERnVsxa5kJHkSgrpE6M4O58/Q2jTvJPoL9PVt/tBmDj
T4vHd/q6BtN6yplR+dkmrbPcO9J6uMD/Uzna33GREkvN8xqBn1DNhey2dopa6v4MRiFsS17UpRon
wocKpsTi1yC1CiOkh1aW28KmcnrbivVZ7HEKEFGsU91ppNf0/bKh3PUhv8Wq+gfqAkz7qoxEW93m
Zl6TIYvMj4jG7voe8PRJBMBFwIAZi9lsXD8FQEQcqbznLUSnyvFc/w4nqW1eDfAAwqXK7r6UgF28
E8BJGzudsVUpjjqWrhmia8PmSY1eqlbYhYf1Pp/ITWV2kt03sZ2pKoFzgEHFTi24BU4cJM2IbOWG
a6Ycs2yo3lHP+e6HFpGrq6gbMPYBnSSGQW1sbnHcRCJSPuvAC2D0Ry5UWLBGFw0fG4NQaO5lZNSt
UEXbS+fDeMmXV1s2AfLE+yyVpoTPaBhuRxIGK/shmNpTvJayncglSL8S1oqlb6Mo0GvNli590X+a
AX+1kuV074vvhahXCY4RIHewSIWNWbIm9s16jniEHDG7VDZ7RdokAK3vRuIC+zUhdmuzbbbFSyDw
eBCXNQpGdVGBDizKq0Xe9D4Ua7oxuupxfzMoU0FdSLZdaOML5/MU4pcPYUVTbjqJAuIddf1ZtVrf
oqQOrXqxRUY2TYUf6CNFyIzWJxqtBQET02Ww6FcrcR/7v3dP2vLsucsD6TRDiSydjrBNLgANfxBC
6SCO8VbFIs5DIMulSOrbJ3tE7J+PzHrmvW/kuNFr2c9NikRK/1zeJofEGug2i+CsZ83t5TFLC+4G
zAJ1Z+J3MvIRIQdIJA7SMVadrJV7HBvcrMFJ+X7ciGK4wTKeHhjz+m9h5u07dNrfGUORvVd6rjlZ
K6eoFD6F0u2JoZcFWzfl3wYXhV30mn5flwLuYPZgII6kD8WNfpGpoopeJOeuRN8bbMi1KaqFeYgi
p2xv7oD66NOyMZeMpBcKCQxXrMw15tSFWVgRti02XpRlR7MFdxcFeWACpwl3rk3UmtkabIlRdm/O
U4ESFeZPxZ12CCKKBsRgk975/xgMubj5I/elUblqSiKJnSRjKj/SSFz79VT5HPFpMus1G8R++SX2
T/+nNrEb9PiOEpaAL+TJ1yVYRY7P6ED+uVfYSJ1uO9UHLx/M+MV5uR6IdCI8kumpAwYxnSOrjLHc
zF7mEIT63YJaEWFEPUj/dkHurccq7jFUpUQpoHAkx+NwWyLuSsZCSnZWW8BHeD6etH80HhYFoYGi
fsPIx3Xpw4ypSefDjgJCaoOx1CQdUwiTEO/fySififxZ8tGYoX6ZUDqEsGCjaxiERHPo4GCYKGOw
mfHrnRMwUVw9MgN2EAhm3zb5KPP/Hpqgodla8KuWctxASXM4tNLY/HYXTV7FG8cU1zSWYzpRh4Z/
XY+NMFs7llBcM00L9iUKBnLjL/zvHYnPzXqLovN2APn2A8mEue9z8lrWhAigexWaCTXZeHJfDuxd
+WdaN05Ntdy/Zj86OWS3Ly8a9JP1C1t0k0rEgQ7o745VCSvF+k4JUrKjsUA/jMJ+ljX/uGb9ukOM
YihLBOXkdoCpjvqjdN41lWnVubqzYhAWZHZY/DEYwPFehVqGrf4WfYGhxSYuiKOc8KzQ0WuB03ow
ntuU0Wj/5jwEr8HN6JEjPE0LM7HoAjEDUcuKJPhCqNNvbki/BP8VQeKij7tgEjro7/asS2ocrsXh
29OlkxeY1LywbzY4nZJaEiLmhtoMKtCYWr7yYgK+wa8U6UVcsfapR3EuGRAVI7b/d3LP/nL4rdyo
j2IUCb7CD7gDh5iXBcrT5x6fcMak1T7dDm8JWDIJwWJbzQhSeIs5vjGLdgXfkFcMHuH54s7b2fOD
i/UKELX3ht5lkM6fANSlZgMqRNRqqktj9gTzQa8Dn5EzeMtCkdA1hbvKiJ6xqQGhpRD7UdhWvi5J
QwP9J3kON93gmWFj3v2NccPtsYtguMQT1qBm3MoUx+QOxVHA2c5XE3pkz7vBRPtn0B6MbO2tRY8p
fXXA8YLxdx+Ot/eVZ2g8Gypyqturb2w7cw28OMAB6a3/jXPr0/fadlmIhJ83DMEahvEFNTTmuyc8
/rsW715HS0Nj+EE5PlJBMNEAeHFjW0+TI89L9Z1x4+rqNlijZqCqyVFMvuPmj371fFZX/rbbCflf
XB3+mkh662to65Q5ZwWp6tDxNYhyZHnzWgzmrCaPWE7iPEghiTMYLvX1Y8iIpuJNirzwin5XaNxQ
KQGQNbTIcMyTmgKzmzdHqtL1TEc09kPb2HF1Zm4zTH/5h/PCvH+1A089Twu73+Z5w0IlPRQ3q3Zy
4cTSj/zXjNwnCz7IMBSvxgr9OTJBbwYa1rJ3TrLL85Fws6nUU/ckmZFb25ffx7bz8CacbkRsL+zJ
gfaokkhAAsp+ujlNutlirajLzYdaJ920X00KaHmSorNhAVFIgwPFMRGC3PXu4RA4ZXt5+Gz5LliA
rSnw/Ht6Fd5kQboOE2nd3aRhvbAD8k5A/U6xAAhzDM3u1Nyh7jg2YSItD0SS4Ea/2aBWFn42+5Yr
AUS3vWewL1fjKDLTbN1zvHhitPdypbxAbxDyhrIQU/U3ByNYg9X5CnZAD+HyOMnpvwutp+715y3L
a0tp9ApVfTuqIWMtnjvFDmYsqKDw+x2v/fjBw6bKieVzq+qgPoQv4xvtujTr9jGi18FHFRT5qmYR
/G8tuil0LReF2XKsh7Hr6T0EuT0kdsRsxUPrTopeimlmUFX5XWOojiBftD5JCmiMxQVgDFagkagH
uKJX+NYSNOPNXFNZ86UMFXODmnLtjtpZmBzuVnQ4IEGY6IfKa6fH2HF0B5s/kOYm4z+4R28Pq22h
32zT9s2nX6Z+i1ay7dn7AXPr2Y4+6sJBkhRYOUE6vZkivstKhpQRG/ZBynzSSUmY2sP2Fd6ArBN5
D0jP/YnQ0WLzUm5mSR4BMOhnq/pGfsrDjycvGfDCkJENZOLlCuKxI6yDIIS2MwSpYyi2PTdxvbha
K4Wv14Dcg67LG6MQlQGTZMDlnY+htB/Y1DnEppZnccqqGcrOpPnK3wd1c/UaLUrjAaP77ExwIOQA
DdTSN4jIFRLsFD5O7rYwg689kuW6rlIEVYgKrM7yKbuY9qI+gM8CC36d5nqmK5kyMjee11IRlT9M
OULawq/Vu0jOYCfoeH0GRrGKCcXRTI8yZA8fmpQASbhy6jRqaaj8ehmMphVuQVfQB7qJ3WfCZAfL
1Ak9JoXAnaETiWvn5LLhFU8pAv4T3SX6w7xQtCGlRKzwwmkYK0rRXDLlTfvRprFsVzIApJTq2Hyh
qg+15Sq3Vhi/BClRaYEqYSIC1/WzQHXQWLo4FHgchBOvFn+vHajMj0aRh4ptRduP6S+Yx1PlYq/2
TEOR6dNm7r0hFnZ3BRe8xsovkTfYdkINkRZbJEabeYRjTDKc4PKGZXVRZRGJA4sZeawuYXGT1SKv
SPVywAkT9im3jVg+cXVBYOC/Or4mUxTyP/C2pN9TDiTO/Gl9khS7c7IjRdpYlPYwyoR1cIeNXTb1
toAM7iGS2xn9LEFq/JxGxF2QcWNrqYhZRYv6MVXBRjGnam0psScl/Zu9mZO8FJhN5V06+92ct7T0
R7zIZrVq6Kr6bA+l2uOt5qbJmntkXwDs6cq18aqYfBlXTv/mVTNCOI0udPX9/vRKsbzzSu17gLAJ
EVxJajeqStL6zlaXr6/V7PKV3x6FYN82YjyGY/Z7tAfzV1SOq7U6WeTIJH1IJVLSykL25eo5A/HV
ourcoA4ScFiUFQmuz69q9wi/sMYzU689ncaiVB5cw67ikCYpX2cjOKiXM0HclO/rCaRUae5/IxB5
LSzhMEEBVcUNIscBvynCDijW+6pWP1PGDYFDAjHGkH6EElhWqWHx64GT8NfV/+8+6JjbCELG28ZS
uLVU+ATqabt5rLEmQPwbsRSKpBsU2FeG2PMd/VbjnDKBXOiX4wiPtRL3x8Gek1pEYHusNYYOlwp1
ySLIfKIMKhF4SOR7FJd9/D52NpUYwsYANlcgL4WuuPDYQNYSkg665Q/cJ7jd/SquJM8rmAdQMStJ
HxzPh0/upcSvkXwWIuEqQxz/lwYH57j0i7+DRy4OzVBZgb2F0lQkjGOfVo3zQmFONlP4x8+YHIv9
Td0MFjs1syn0Pd71flxp6Xo8WXQaMYJ1GBA43u9XNnC/7z8xRnS0TphkIRUBv/kgUPSYuELzbboU
/wuRVqHtUAGQdOXiHF3kvTPl95OLWbS9KdjWMd7u6etkK0+E/3c+IZkI6mk68yvX+w+WA2oMjwn1
66P0GeE544VtkdikRS+9O1++YsOaWS7wu/W9+yQ8wkeC3Lw0eUzAgD6i78cBJaDG9Du9Ii/trOv0
E5lc1vquC1kHEWhxOw5adeZMvkXQFrZMSj9uta1lMZrT5MiRr6r+iIzyrflChNSsu5eGJrFfD23e
7WZPMq52MxI1W7mtP0kwQoX1QZgo61zsQOFxhqNrPG2ASB8E9tXe+5sme28/we96ABs5mzu+h+QA
g9VZSQYFiOZfgVvNErabya66POsuS4zr66hIV1M3HhOKwXI0vz8VAhWFgW5gjzU8OATrfI/8Tduh
UNZyZBJ25imNshVeT9ZlqhPVDpIguW4rRFHF9OVC91DBm844SbRbApby8pecvnWPxnf+PRafkXj3
Gop8rgb2Gtw/wj8sP2+qiRTjGXrLrm7eHcJ673VJHIPX1iiovZLa8Z88rJBXkP4/fHs/7LhsAP57
A/Kr3Rkg85LhPECkrfTUaiX9pm9tfsJMyPf+dvtZr2hKcmByaW3s7OPtr0DrtqesDAxt0bXRJzmH
pLJBb2/H6dnCMCCVWG/us6MV7HJ1v562fOC+6JUk2nhgvncOxetZUUqmyI/glRmmqK5o9DVW4c2p
SE956jIbwGrYAdNyyGmKUWfcmK4zfDJo+6gg5vZMA1NPHbkmV0WblLSqNvWnUdIEjZTHANoKI9Ml
4mndfIFuFtp3zUomy0RbPmEvTk3CcD9QMzdqlOroBOzx0MCitgnb0njG3fNxZF7k2FkKZQbMoHzJ
pMOnxqWuNTEPZ+7e5Km7OsJLjDGz2v5e4B2a0CtiW+kiMyHZpnelLxLQAcfLYx950aswZ6RW7QnU
kEBxdclWJLxmDknM2mH+kcMsftxModK4w+8627d90WJoCB+3uMIKJZlE5qOwsbesSIT+JXN4GszM
H0EpG8Jk7Voc9gzvqvErUxD7YrUjYho8UNxSVnGMcwRn1GLiHdaqN/XWM8KIQRsJVt9/ief60lac
EQeu82Tmpi1s6QHPWvrCguIMjpVX/qMIelDvFK1T5TdT1xw3997gpOAsmu7Y2u+PwFcMva5LEGi0
4chFTObOj0J9SgCy+sK1wETCFPNLp30gxHH1ksXmqYr2HAMu0KCbsVaE4BnX2gj1PQNGZTkUGq2b
n7LSXNSmJMOPsGrBELLtdIhNVpZmshfbid1+cnBANx4Eboi8qLXFD/HZow1WGhon/G+zdeYvgnyR
e5EDB7ffZa8HIaZgOCsBGqCj/8UO4EiJ6Y9lXqP2CSzjZ+MphrYLFrygEp/5oqgPnVn2yK35TY9h
mEKA9H6y9fVwYClPwkwB7vIGQ9ykNyppIxDFvhPT+N2dYMTBPio78nnXNVcuHPIWORP53bmXPpCy
XnMLUtWdvJZmF9nuUeHgbIIPPJYjSPh0AUJ8gFmUl6keIfSC6Gtf1zYlwlLoz45bEUmvyMB16oPB
XFSCovykiPD5OWHARAmSQG/nJaseoZR0yy/e7d1mZvWci/F3jWYzgVf/xSg0JsrXrszVSNKdxybL
DaJbqPWP8faz9+7/j73s5RI0wFZ0KqO6dZTf5ZJRL2KvUCpFmdeOXJ+YhtkMh78t9Ymm/oPZ/6MY
wkwST/bS26RWWGNoZvJDenKCad6GMyjkDWEdo3WNpqVaGaCRi9QZioY+8z6fQzxelxhYwer9q3X8
yV9epmhX8skfuh67k2lG1Cw4eoWydfJ6qM1dcwn+o9ooRjsYhecAkVZQ3eVHV1GOoyJ2FZo5SWH2
TE2J7LGTT7VCnCCyR6QVFeDYL4DoulADBSxB8shg6UIUMD0NWvUIKHHwcO+KH7EG5CP9NjSzq498
FKPJNLqQ/kLRP+QUJnWKNAmogfycXqqeSNr1Z4maCv5zUTwcsska7Obo5muz10797v/btVBFI78+
QDc4/GqXLSL7kfcorq2yXCvH7xK6b/Png+5ETuWKhl6oyLtaskBYHP79tjN0zpObiNojcTifZ6et
0GAW+Q2qDBRQdLOmj3P0izk+8rMsJ4KLzf3zyF70+r8staJoVW15GqXg2SjA2WhVC6bpbc/34AwV
dpMGvMJ5DfvRfpXYvtg5w/qXubimg+tRsHgB6D9Nunm0I1sJrR7w+Z0lPSkvnMKT9ne7u9rsuhbJ
iNH7h45xZ19Q2ES8DkPnSVz/im95N6L827w8BrPr2Y2BAOVlyzWfJQ7He8wYUpk9He2pQChOk/Id
k3/amti3CaU67YBnyw/7novskkl4yxoSTX7OJAD4RoaAvJwnVWXPFMyXfFfom9HlxZJGKEm2Bm0L
YWH5y/q/hFvKxM6XViSnEcv2P7lDdm28FDoH2ZIyDghBn8BLtlaqzsJK4vMZK6V8lTJ31n2sJHOo
5cixqJ+eMVR0O/gjCN8RhvzRZgcPzDD+SRAnPhHLK+LwdXCV9j0vPLt7opwIbRnh7bMRc2Jmlc4v
3hlj3JgAPsET5sMWuMzeXvWoKng/076jkvuAkzliiEFoXC790fPf9G0Qj8PYpfbSf0+fwjLkri5v
cRfHjrhThN/Ykgu6B2tFsjRmtna/r/DpW6RbK9viAjG4SRBa5s68ZUMtfGHYjyWqPCmU8XkDO/VK
vchjPjP+GaQYRYxKY9retJSpvlgp4sdE64nFTMYw6SmVC5NdCjMjS23j88FGhMzBwkSUotbfpL0l
p0v0TDP+V9ZGr+xQaab8RPKMnsbCmqjJA+9f9gBqapQU0WghgZrRjqwmG8FBS7lTHxsSy4gcgunR
PVBfOm+rWqnrQuGQPwXr0LmN3+dxrty1mX67BhSH8515Yot97viBxIp10q74g5ld/QeUjPNTTJIy
luRaG0e279xtREO6Ul0LDpMGIryu263cOV4g5Us9jXc6k/dw2q+gbgeUwj0X3tkX6UZBXbuujGyk
SYT7amc9sNtvzvCrNbTitjMtDv5Yn06z87KtJIbS1E5Qw4PiG7tAuU4B1lwuCRhi/Ek/QHhqFGdW
PH9WQk+OwT0zXOat6MJfI4DVut+hGVmpPSfjLpA/5jJmsHr3DP9n0UGRXG9pwDxAd4rbQ4jexi5q
X/pv7KrlgsxXg4Bh2AZwq+CQmALkz2kLyvbAEbYlBWvbpJBF7zxfTXWQvQdWCTbP75c6L0dWAG8q
qs6LhuGaeIQXdOAmSUvfnQiQI4bUII6hm41OxiJotu0JSK9p+xVCkpQFP2g7ddeIRFi8FrSxerBE
7PeZ9MFxGEaoBUGxsx3JPsqPONL0ARx7No/x/3SmPNAfqhcYMBh0KeTrJ80HJS0Kmf1nHWcOuAHf
Qg77NuQxc0BV2wbdMrxOeywSsQeuscJOMMSfEioepbPoRS2eIAIVUzhW4YU2omLn6PrlaSY2jtQg
FEj8Um+ZKdseZEkNw2U/rRj2OXkHajq18gn233TpMqXD2Tp4nERS503uB9WOk2SGgGXz+7kDchVa
KtAzvyLXCj987caTuPZTJ+Iiae7cxqfyCZWxPag7asSQl/MveMjZjAcZqv/UqbaMKNfyt0XOkD+K
7J/z9KHw62HwQGo5Pu3gkcMnAOI9jed0aa+5mWaOCYkMhqIM9B8qnymQeBetN7TEiQJd10HWQv44
KEAJstdWWwtp9FnSnFKyl+5fi0ZBPg6BqUC6h3iOvn3Lew8qazNTbhgKTfxOm1vP0jvrfxhpRLWr
6WpbO/+gJXZ1pfrPoCbSrD0gsBS5mPETnPYjis916zDA+oMT0GDKl7BfPOYQVs3KlxaJqNCMC3jO
mnKaQowbJLRpeZave6/ahjvkovVbxjqpYTYKr1KmnF0UCxt5dnS/9M9CUaq6VkRs9mVsLB8BOAjl
EYf9WeymRTXViOd4S7DEqe8vZeYOF0NDMqtW++ujLx0SxEInAwicngNaolgWoqHRuyje3eTjsdkn
jPyxiO1DOMS8YZDMYBgpD2SAC2wUFnjPCw6FlFDkSmVgcMYRaXrPAPuXaiJiBuKg6gnlzgjwpxYo
iC8yuDPEdZN5WpKa7XZybTS3YBqAc5g7JiwSN6M/Yx3McafyoZsqONn7V9Or/K7lruHWa0ccWvrI
1lSlWYCYOd/v5knDWtPJsyAjlGDdd8fepp/fOPFXsJD8uzXlXQAM4BgCPbSoDiprPdENG0pmFGgk
bp51r4jqYhPEquJtLTEuGkgEHC6/6Xzs+WAE0F517HI3rokjrtlthhbBHefu4hK3fbfOjPqzYg/e
j04pmv+JnUykjhykRKerZmra3Bi6qTVPJjdBDqIjCLWHW263haCYILaNoAwX/enVMg1+n547bfSU
2JA8CcaFHF95c+nGQMdt4D7LK2Td/sqVgMo4NDdfKzAT+UPFbP+vtJBdzlQMfa3EhhZxNwHu4hLv
XQoByQakSCGcu1mzNIxEzhQpkVPwuw9plfjidpm4xwEKoUdj8UBVJ/W9weeDmpxRSzA4yTXU/XSc
pJW3ruW1xe+EvL6c+10UEuNCFCyGwhcs3LwcZsr8JGyxNu4L4+t13IL6LU09hXy2hFMhjzV2xrgo
6GHqqFDM20gJansfeYV3OKndVUBWoilNB2DXWLpDUd/bRdVGpQmmsDcGBdGyNMIXYj+IppujijL4
xiBWL3YgPYdsiHt8f+PwEzQCxaQN63Cylny8lkMAOvNWPfhXXxaKWKUxdtUgVUA/W4pBu7byYcZK
OSQ3Flp5dgSavKF7uqEAcFQ2ynYEpSyTEcmTWQ6lUAC8ppe6ZHhsPvQgIPS42Mut+E/a/w2wvU5D
/qpCSbNMdOK55qLQZMlefRvirdsT8Eu3i4Sq/VmjzUlqOy2asVc8jq+nWt09LsKBDCq+WEwFDMaP
+dX51MweLrTJBHYhiHEiJ/UkC6zDxWDCfsSCo69Q9v4gnU5CCDAcVjA/nIMVAKtssb5EoIJu+rmm
h3/IF1FhOxyWUsmYrRrhumZ7Ln5c4LOEE2da0KeeaScYdH+JzAPs6lul2FVnqtSUwoKdf1srLZrA
f8MZ2R+kO7LWmslHLanruJcpEsxuFRYjbtTJdLM9UxabowM1DPkzEhGEigTt82uFPhsxstgjSnz9
pQT95WPoAvnkAgtYp8hATf55eRRA0pEuOUm9oIJ6bfdUmsuvtcenlUYMYCE7+gBa8Zu3Trs5J/Ji
mKMADG2zkQA8jYf7qLHl50qWfpYHEZ8fOLqSLE8ZgzcsoeA+/H34v499wGoU077aJvPGVSIXJjxs
/uLcQCgLw3aoqhjKpE9jE/sba8Ku2SZyh6ynsu/r3SOcZRf0xA8Xen0vZeCPMEV1dbDuhRoJvhLM
wGZ5gwvpP5/vh/Ju1qp5p5dJUy2tYdrGrD4NwQOc1gPr0rFcxlYRiNWXtb01AxLlafyBmSNELZFy
wOL11Po7dzwKNSCu5TiuN+yjVen0tMkDh4bG5yY4Xi169fmaFhU71fmr1M1sIZpnITMRVsIhsbGs
ChW9KtOhnD/MB3r8oFUcGZJ9waWTLcpqJ8PnI7gnJS6KPtHaUJsJUgfPpiBXB57A8wMLbvt6RtRY
z5t2TpJuQcVquapmJypNaci6R0Hx32w5qtR0TFR2+CdoQVuyCOgv2BiJmNf1EG7hRIEHjxPeBB+2
LdRQZ7ggDwLk8d1Gfke1LvMIzv1L9/jNJDMPuKE/EnMqAiOlQKL+qN/aSPQ15xGl2GAyDHwx1iRz
367Jfmoesl5L6Oeq4MOgqDMUIMbYjxo3wc6Fjt1E2lADO/qpMsbLzhZJ0631CTH8SjGnYfx2mjBL
bIwol7f0QutqGVG9JMrImA4gh8c5CyCzjaFE6+L7AjzbytRVFHFZL5pMWAWSaapHd60DbBNm1zXc
N87v/DPF0DrsWgfij/mSZBcPtntaghvBEHqN7MS3gq9WcIk7NQ1zqIXBFBS02OFbe5XRmuQGvhZF
UvmvDK8b9t2GSevhNSHlkvGxe1EZi1M0L4EXweqlxJZqXpYEErwWxcD00pkkIslgt94OJkKtMhlK
UCcXHvp2buBSgr5UZCRstba+eymtP/rFimMjrZWgeEPZV7lcdQag59q/lv7DFsiWjOhOoDzFsbKh
r9GIO/LhKz6/tENdyBEQRiK8SPWWyrRuTzMjuDk+4MtqfwSlyOH1Y3XqAi3F3NdsMZ2ya9QDdE5R
tZdC/ibcYU+GOnX/cmtf8H6/wcWC+Ln2qK6AwAc4L5qyS3SzNiukiAaTLRcYYki79RMGr2kHJgbT
f9BwooAUn9axfcSmtT9lIVm6EXBrNUPtfxI/HuvrA72WMlP7KWYqnuKJkeVqoK3T29dYvNs9A7sJ
6uVx2IzsxdIRFPBt35X6Jg4JIy1B1n9p9J0GerDYlOrQKzTTuyohAdUTrZeJapZhJEMKKzR1E3UH
5LuWHc4D8edZ4P27We0d+EGRt1LpYRiDp5gPH3wPxyBhWVosat9s0hC+6zYaWRL27FWV8j8Z1pZ/
xu9FYIAnZuem5ExQCOafMcaIBy5ShmRuOqT/5oB3WnbfFe1OKka9hytm1VqqD3wQEdUYH9L9mE8V
ln01ZnKFxcUp0NLJVaBnYqb1PXxkknJ3umzlwJMqE7keqdrtPvCx740O19olMdsMtq/APYUsIHgd
HKh7sgHoj/UsEqghx3JIZ3JTK3DlwuJFBnBcLCZTySo/NrQw+r2q1r2a4fedNcwZQSi9KFVFTZ5V
Nej7L+T3p+tRAk6riGSRD5GpKIR0Z0/WsCXtsJc6d9dIZydl8umV8JKV6fhIDWaproKs0yT7179v
LUiPWB10csb29u1VJnpJCfFzFMN6NRnKGXsNHJpaumz9cgiAuOY8eoJ+rHEgDV/x7synblkIAjNW
S20wMaLTWX6F53SngPncn2dqUQmtw0bWnFLFmpDYJMmgIQ4COPQTBLJ4JSNGqLFCV+bB6r6r11EO
kUMOdEQj93L6pfBSg2uxj6n9wj7CVW1vvYVFOhNn8hwA7XT4rTJSVsUtd5IVLrntnLooPEeg4NXv
jdzkpciLNDDw1zs53gO6z11bayIBEpdsyHjKf7Ieav8cymVi0k0ToavpjP52iPLjX3i6mbly3NzI
G0TE9GOjXdeS0CIX7RJzYBC0XSFCLU7GncQXWuH40nEgm0+mYZx8pKHR4cleyl30BBJQBp9p+Ulq
tqWWLFQ0wzVnh9NFaSLFoF+UDJ3xFXAzuhElrIjQuSqABxT3BiDDpGZ1EQuuhEMZOZZjlB0XKQav
CSMV6xEhsIGI2pN00XvTdRwF/TK4ESwWXiDUs9lSwzy7AkPYl79n5chEJGznWbfWDMzXyQ5fLmr3
KiRQVm8e5/nbcFaP4qRbfRzzgeIFvMF/1oQj1+XE9+lebX/wpyF9ZrMBWYEoGHG4PqIT2Yq0QQU3
VfodFGqB+5IkXySQSAiEU8EjqzA499wvmDMIi8NCjg5k16O+h+z1lrz7T0naAVilWyL5R29c1S/V
ckZeMm3MCdqq3OmR8GQoR2ENcwK3iMXS0AmzRGXKFEDQUz0f+7P8dqHMGBsa8lRLXUHWNQR/3c+5
Gst2M2lDDCKFRUFsij05VHoGCZtomz8bGhJL52v2tQwBd6LwfEM3kkDJgn/Ve1r8ug6I3Tl84Tsv
7ats2JoPVj7OdpvnfU+U2o6eECnsf8noScXbmNEevCpjS8sIm8sZRxytuNJXvHS64KTKPAPRZxTH
/QPfTNhQDoNU4alEwGLB43BAnyVQTtKnL3gx7CTNf6lRLsHhOlcpfJFQdiJoKSA/3q5BhI2HBzRA
2UcDxfPffZmqwqCSHYlrekYTZ9qGFvAbgjzkEN+P1z21Hhau+xnuKT4rTZ994MClrvUcKi3V1Xsu
ePiBPdic522XB1q+T+PYJpveKsaH2ZH1r6ebpacUWLZJZV2cztDKo0InQTQZUzWOrhggWetaNgk1
wswo6dJl5Lji39ZRqCKe+xZ5AYBelJJZVEmvSu9N9CMtimBMPffQBvcunRbEHX68Z9r1lH4gGtev
dXXf4asZCTlEKW9uS47TGCBGnykB/+SHeAo4n9VYaiJ7x9KY2Zxk++vny8/Hmk8epOPPx+MKztE4
r2ceAaucKO61M/2r47upXsZMjsexUGAgQ59ZP8UG9ZlNNy3kYGZs0f8ry39X4mzeF5jg1lNWxbT4
0MGee+VzakshdLtax022u3/sg9L/9phZEuyAi7v36UXDnt0b1jk7uPlWBZjKO/joHoWHmsIwLTvC
3E/L2JjMT/99xjpqFiGp1cYVhFApbU4zQgNbjJlBC88nvPgW0cwK9ifAeFSg4njaUkfR7drF8vEn
WmjQwNhCy9mfP3LLoST4bfB6/XAfH2QkN8hHyWHINY4Yw95Q3yC7FnFcyr1iZRtjMrGjodjh9t1q
Br8HMg72bl5mRiS+vf0jZm0bLGTHNNg+nKqaMAk4C6QB/9Jhv59qP0NIE2SsoUDUi2Q4sfMTyvcx
Q4YJ4e/ETyk3V1vOtPK0oiD60SKX5muQSNIW2ZRzcrHGYysKblJXmQtWrczDgzaD9OMswkGFTjag
QEduNusrduUOnTJfi0XV6OqoLX5V+mdzLtUpxDl6Af5/GhPfhNjSoxo4+nPBXxWtvHSLW7Hd2w9B
1xbNb80jxet2buRC5jSdY4gPf6yTFitjcTtwZN6C35e6BzJUF7H0TUenvOGcw47ku9bat46H7LDP
z39wtTdreHK7bUQMyhOLpuk535bQuLIQXFGmHhbWsW9E/hO5LF+1PVeAJbAfUO+3WMUIluSJKx+i
W3th7MYSchtxOXvvyenUBKKyo6LtX2LUmtjK7yp0ylmBIrDYU6rcaRWmvUzV0ovQzEGrBFDjPT6b
ObFqzNbOBAFR1egxDnSMXK3eUlcC6FToRhQgXkIZugDPHVJI7e3PxlUoGSnlxccEWF32h/gNEcCe
b/4nXtDgiDnWDZ/TuhsOVtK7zRhJ5ShJeBO9A3yr4PuJSPGsw21/T8ptJvHE4egiBw2e2fATAaon
iwMmwYNcWio9hzHAzbkYUvWa+Qx7dStsOBTFll7Y60T7UsXEkivslC7HTwudzzTpDpH8IPw/o00o
w+qiUexd6Js9jbnupjzuzPsZvKN+B30946P7FfDXejyhsFLKUK5IPWdmqe6bIBOqeaqKb3VnD5xM
N0iaiEtN60N4L9otfjdTMF6zqfbdxTglb/YGYt4wVZjIZ4ZwLHFU3ebRQHpRKMkcJKLdnWI5aM8p
ey1kqXpNeI9ulVlobOIzcJkLRK17PFRxaZs7FL0ri6Z+awWDG4oSZZyviHCWKAyPADOdkL3PIIN8
LroBEn0TjLTFmWp4lpHFHY9Yjkt7VLBHfre2G/hghR2FbPMDZECOOuKCBSiwSQ8JbMaZoUaPtUWA
TCt1lW7doNi9eX4FxOso7gQusYOH4ZwK2HsMG4hz/5rvVQA8k8fECodAempodZv159NZ4iEJydnO
+lmW/IL7ZdDlnxo1NFkxgiAekHrHQt8JRsXZzGTcpuFVLLCL/flkrCBDuVNj6NL6PnmBPZYMkelT
Yhp85UkfxqRvWOlXZSjI+bqMsQkBpgUFB2CDdIEJZI5By3OrTOooU2UIgGr+SxLWqIIgvANOfO68
gpbyAIw+mjUJS+P5EyDpokGQswKz/yQ7Z7YpUKRlUOrxjsCIPNZAZKjZFimsbgEuyWM22b03BSm2
tOaGtmVq+1iAUYu54LGIhdzv0O5O6gb/zwvnsuJeeoc4/oVG0PUT7NZaHfRz0DwpNLE4lKXvvcgO
AWeCfcENpeARm38nDrGzf2yHnCoDo8nAZ+tflNpVAzCMgF9G8zfDz2MJkt48oSQUs3pJ8LbVvpev
peWSo730+iqZ6zWy4Uep0yeMt85EB5qzX/TAw7wib2ush6gBZ9GUfeMR4EAWBWLrAO7Kp82bf86Y
ap0E7/ca9JNMT3iFEhdmA76VrzvuZzmhrX0E+SI/wcmNzpqNU6RKHMoJxJN1FdN1iPutmwBYKyHo
X4m+uSAtjocpT1nUCWjgQ5IBbEnXijV1Jlq+7PvvSmO5zxhftoxU0MM43WXGN5EKqM7q1W4jToVd
dn5j8p19mX6dpbpZjC5iBWInVtpUSAZFvqPRoVMe1BugP8UmkW6ISYUu7Sd5kt4Sr57TZDlr5kOS
f8tazG3cmNqHdYiULSN8es5S5AbPPJbFCe//tfMdNZRlFoqPc/oyvSGyq1wrBYLrLRLHmJp0sPuk
NyHuln60shevFNyrP05bZGCcHiE/MeNRCFNlZCG2r2GJrHLEA0prDHoDbG3hA4z/GViP9ZhtUnh7
8JXSDum1+oIuylT8Qp9nbAAoiYzvxjiGduGYCZ2wO2fBCrji+6xlfih92sOT6BaU8Xxvioc/WJZU
K3vaUrjorWxFkIsHuCp2ACzvm1SPxS+TmRpfDC0X6sr/tlWMFrxvH0We9bdZgId2t/IOxae8RH25
zsI90w1A9v2ICkBUK0yo0luOAPH0SXwqc6yJFF/ax/W0ojQ9ihPhE44e56xrAbqIDZ0x9gLphXJP
hBfr9K0j95wCNfK73MescZzCXtWSoz9xstt/AXARmAW/EfL4lZdc+Gm0e2TK49mttHV+/+6qCeRV
8CuA3sLH7CqcfCb+N5R18Mgcp53ioFo2uId3N2ALU5/MtGhGQOx0bOmOAgxI8+H5n61Co/GVc2qU
2nwtDutHrwtyHjx4J4VpLWY6qpykQAkh6txYIfMBAiti8Ddr2zNfOumBPmUKLLwFBZJLkf/wgYBh
9GK7tL3cXTysmMabvHdOTTnUqUERrf55JQ7gLFiXt66X1Rmmc7uTnPUcsZZ7SIppTFXzJrqmlCCP
nAVfRv8IgbJpCkWG/6sy27NUC9QkoIj8lu1r8RmtV4EaXrLh3BZgdyRMTQggnMAmhXNp4qurn3eP
2Q5+Z8ZD6YvnepfPJ2DNxZClaTlmO50v4XZI5ASQ71+yOdkXfOT34jbgkYyGiYAZ0R/GTOlXNcjT
o35Vyc85PhQXBQto64V/BNAHpia0uTlYYdMxscdswPMHXIX7V4lRadcC9aY6myfqRfKHE+IwYJqT
7YfsNzNdUR50FcPpY46g4Az1U3QxB26akR63OB27n5i+bK8Ge+StXck6+RhLT5k2NEaZRhTPc+OH
v61InF4hvf1cIXofQ24x6vCOYUAZ9SMZOFofpDeH9JfKFN3dh0L3tgbqgoaE3XS203Ig66P5Q5dX
z+SB7lZvuWmQ+WJNL3PltgQZrXLA40x2XpNQOhvqy9O4OBX7giAtS2U3YFF56luyA77oy+c+ta3U
AY3g1HDFjVSLjDKxgCAowymegDKOuTQ3fS/prGIMaVWViHKyNcTHeehp03YENlHcXp4uUsAsz3VW
1uyI6BRg6HvUnh00LIgL8GV240kh0Ls4mBg0g8vpLN7pHJbvLQrB6oUhuPuwNw7oDYLYrJwl4Udy
uQvCsn9WeSQ6lloWgIZJxAlEpXd4kaSRGlUU4OQJYqPCnQayZycKHddANjle3uoqy6epIgrGm76f
dZVN0iR2v+dtIZoTzLd1gA7gWw/Hnh/PqJ0IA0k150u2Vy+xi4X9aZxtNo6GWlH7s4vaLnq2AhXU
Pzz5wlswbxDknFf/ysUxZF+Bs6e7vxYhjEORXxdMmzwVaeOh4LfebUBNvYOkchm69t4Ykb81l6l8
grvz4ddLLO0cjRbAimoa87EiNHSjnFXqR2N9VBqOBsLi389uDKMBgi4GWyfEgnhhvopOaBJMTBJS
is8ySehT/Ku45J8E0r7fnSLfza83aBIX0oG9WGxZZWbFZdjbUqgx4MATL/GvRxD0B2DxZkaVhBOk
2YP1T99WF3nPAIgUQpavVGQ6jL3tAyYh2NGziLbnXja6NcNS9E0cwH8tLxiMi1kiKZeC0IUfxAld
gFvp4Clvdtaz5RMI4txke3LLtitevRfn3GbE3Kjcbg0SIS4VKKFTxelbHH4DBYpCKpvk8Tv+IApF
5Dc6O8blxbhPRCxdtFQqzDYQpfGgMu5lBj04DrV0YWBx9VSDOYMJXbpacCkFxJ7w74uevlQFMAeU
r3NDRLRQ5t32BzxP8WjQc9c0S1lwGP/XN0cndSZzEmTZCNItTPFAK//lCjbJoAQ9JM9sTuyP33kt
7pryut2/PzHmY1r31XmBkppCUlHXrfF9my1UGZA3g+ZRO/fzv4bbaXQChTHsGZQJjgXgAHcFB+UJ
/pajSgIp3z1zkEGGADDKPrEhvds3ZPTma5LG7XAQkGx8ReaAJp0i0fQZI+EqM6zYUBHw05SMahTp
PIA4Rv1YHlifVajhtaYadiwl2djltTUgq/xRt/vA57wtb+AbiixfKlFNe6F3W1F7R6HS57Ae/EiH
zu+lLwlPl/iqpqOVWwleB/R+ia3k0JJbz06O40JRu665bv/kv3Zmjh9dOK/u5f7Sh77NWRlp3shD
SUBXbiA0nQHYEV52by7SO1LDeiU+kzjeWn/lb3uKS669naEyjdoNj1shtsfce8GFzLcMmPtmhlVe
isROtn4Q/8QPgRw7yWb6IEhPErluJxf4rSxk8ibvj85UnW+gB8vljT3g+K9ggZqaYANpjFTNgR7m
NQ68irQNLBLYXdN1Z7iWJtErtZJ0G3hBTZdeVT0SunvgYnsal0eqop2cahAIEUnHQQRwhP+g0B24
KC+kGvQKfICHOLood5KQyYgdMz/7Fj0uy+DklZ05kLAAJaohz+j/YqbRbvB+uT9k7Kiuk+w2wirv
DC+FI1x9QxGVHm2rMgbL4qoz3tXkUY7Ex+nlBy2nG3LbpZmSa3OdeRvLwwbbNDAZJLA1td+Qapyt
hc9BDo8uRQJfL10Fcf26FcTY8nb6iTEoW1LNookECWqvoApOQlgIxb/+UHyTkLdOG+Arzk5FWkpY
kOSznlN1O+7xOiFj+jJPVCIxCR/TiEuKeam5tNtX0iSQKGq2X+/HeV1KgjwFIvj9WZiUvsAxF5G4
PfLegXsluvMS0hJ6N1LLj6047FHmDYbfppBPOPRWMUcUMVOgkcYk7WmpVnq5XymCsW1a8rBd8egv
EGk0jPG9ErlVZdGsaZ3RRN81lRjPqoZIbjnUM3G2EfyniULAQD4kQOLEVxzCrJZB1N48BtNLEnih
ulDYPHScRhv0jqHC6pUUN7yTRnz5EBEttMfbahYN1oXTAjkhn/wa/Pylt7cVILY1m/28N7Encryr
BmAvPYDlRRzN5rg6iPuiYFnJ7YDy4saE7PvtUcbyOUEyJdgNO39LA3zT9f8mB1c5btlqLKSLhpjj
1Xk+SrsKYEaq6vVOSe/eBJOE2OWJbMgIzAzx74pxE+uXiqM06LfzFCRE5TGJ5kID0aXtJwEgMLCv
Trik33hcOcp/AmSfd+XRKlMWgID4wFCqy/50BKnELobBJT8wr4egW7TzLcoJm2UywS38hkc7zt/l
NJNRwPB8BN0g7aZH68AP3PEK3hfTsZ7AWiba3welftswhiL5monYHpPfm1tco9Xr5PuGok/JV+UL
yK59gcbTkBkjOuhoJ9qesA6KfM27pzML7yzhc3hW4zBZ8XesFCWwgR/MtGVe/RlZp/xACtGn2RE/
/qJSN3gKe2AdQeTbShZo8rXcHC1qNoNtsrJKqHSvA+/QAijejalh5K/AV8RVK2dB/5Bl6YQm5CKJ
Og1CHxrHQZApyMb9dGCN3SEAPzJ/t/gBgreCPdjDUSo4WCnbEl5eaQGmGHTuG4PpkABAz0md3+fe
41U3hmic4/n7WI+9weh7LNMdEHy4bRn+Db70ztnLxVu3PfPqjv8VqNZExB505vmQ3oYP+aKrmSMW
AHmvo/eRhsOvG49ss/rXiAspWqQtgvqdbZ47cL3kjW1RBJbeYkh3bIdxOdcm1LGc01D1kjIoB9jh
b8iPyagY3tRy+6NZO2iL6ff4u/MOtvd1Jf8M7XVuPoPkUUtWJj7SXecN19o/nKmzQFKjMQROLrO2
nCdqQ8ygogPwSYY58u6yAo+i0zCW+VNNJjTJ9wKBeo3XSkAsLKpOhF6EkfIMxqUDTzQUeqQL/28i
B4KCo0iWKk+Yc0LLNQ8n+r3Czp7jVZreG6Sw5/5XN7J8JAS8ZWZR11mgB4AIpmDj2lon8r8B4Je1
isqmjBCqxN65WXdEt35Ay14nWDbPaOIfzZMAuaRJ4geAW3/t79Ew3OExChneazsFC6WMUyarfyG9
1necdv7GwYUMokaE5nC2abo8illArbVSxZY6QbbNBOzyFpPtoIee46W7tUI+jbEriJ0qS33A1iac
WOB8wpvhsr0pHTWGDCnMLn4csPGKSQvDD4A65G097WbN2fEj5pAoadIXg3UrqioltfeYoKYZcBRr
shNcvVxBlo9LTmXBUbXyOZwGi/4qM58whU34xd/g/CuwE798VZCVELajyoHc8lkmuxk8qzUyfzo+
EpxkERr3+AH5rSpvE4sRhakF7aky8ty85sExsBfMnoB0evRur/N74su1AxiMz8Kef4Vu3P5jq54Z
Xee6LO5lup6QZv33j/bLc0Gg/SzQGvZjEk2M76bGJINDeGRZO7lXDKlMtJgwok4wFFyQXqaxutOs
BW/6WV4xOT+ZeEcWIYlA4XPUPqBDRlOd5rCFUTjw0vfprRGeMugj2ZN4m59q6a8Hl3Pn5x4ZQ9sf
+fH4hyzXv/2YGzw+12v7Lz54owq2AvukCa6U4ORYMP+0EwEDSzO7aHnWeqoGRXgxUiZ0dkoCHwQs
QbkqyUlaGGzk4AQusRpGzGGGos1LTQYzsg9Pkeao6LYhQoq6Q29MdybyYkEZr8IYE3UmJmJdufit
kff6strDIs96a92sAPLm22TgwcIFR4x+f2ImslHaEi1zQji+zmYQnbwfN79oaUq86bMwciUs5yKC
irLn3vnbvKB6Iqd1vfvvcNWkTCp3AfxeoveUxZ2O8JrL7LuI5JYZoplSPrxxrmdcuG/OsKEBNARo
ejx7fG1WAbFbEPT4MLzP4h5z6ZarQy6lQr6rPElR9aR67/cyQICxRm2lL2ztSvnPUmNKdE5z+ptv
MeTxMq6gLdT5OKGTVqcIjWNAz2XjBDp5fEaNbU4lWPefiKK5qSIQN8MhZ6byLQhaW5Mdu9d2E2iv
K/Dk6XoBjvd7MkXp0gYqpHU4nzRlKRDD+zg3gWbzJ2IqpRLCEuKL0RsrmOH46ZNhSWDzH5RwYb3A
v9m9fbYMTUjSRcKvyQhSBuLR01KCZ0ewi+hKKsZDBc+w/ug17Ak6iVB/wTBonWkjUdFONGyqlSyv
ZfIKZjy7Vd2Ut/LRl1fjhmV93B1/y6g63gOF2MqkEcx2N3Sw1hzUBdTuWPWNG+M3Y/5Dl5y1K6as
t6dpyfEXD2NDFOC8ODoyAZXVsJqZK9/ZBzTRpBGFXWZzMuL4uISC30JjwHegWLSwDGNi2Sa8v3hg
C+z1SduXpF3HHxYUhlHv+clEM5XNkZYFmrAXcBAA0IFGoOiJ6bbpB8RPJNQS++Jt8cJxsjEhqANo
WeMqS1fgUd2XnkN5jcdDbrYFv5yRUuV/myaNtx6qzRpKo52BViWVqibClQyE3i3LufPHUPNlkaUH
1f8e5kMBdQEdlAzxrx+6Mq5FTCY4W/NIlFEOcyN0odqe9ZmAunAdPMDG8rf1WZtRSNzV4gTDaChy
DnkkurzsRJow0i0f/en+LdPX4SQmB/GXwiBdlZ0Fjwc1uksmQb3CgroqDEI69rzp4uDFtsY0YdDW
0qvta1fvZVcqMBUuymmsTaxlQnD6y2+RkYm/OS1qpWlAU6kgf/YyLB3EP5BF+i33Mfam+wRRVsqO
YhyPEg0SDjQNDvNTQAtZAfM9qQXb3vnR340+rZ2bw/3K/3Ugb6SUEf6+1u6IYO5GG7tzS/x2yaoE
cVi1RatVhzUTkTIqN5bTbRCDAyPx0/4e8Xlab64Qr/v7LSHzsd0BsxVFh8mRjPGrGGJiaKCNPJ38
m5XzyZiX3qPyG7uj1Bq/z34IOjL9Ffa+wKX+75kQwS3DjSvk2GSxeRM8nUOd4pM0Ltbcyx5baXzC
LUtcKANt4sYr5thgtPszubzCzyIbtXeWxiVZcyAss4FaDTpDG55BL46Hv4TCs+yXi4UwUK8wHm+J
r8rHHoUOWP7qsfVTxtL4l/v0UVD12d0db2kfk17GqDniRN51oWkDNXSsf9n5X3BujJDADSlbJven
LXFVN2WskklxgMftMjeZxiqUPklJShzp5Ecnf21/wHBi1E4WXBRkSY0hX2PHxSrgWPDspU7uXjvs
tr5vnE10vpOLSrtBfCL2KK6w+XQG8r3/FmiT+XyBoMmZ5UXw1yTZx04MF/kUdiSNURTVZhv7Hdfj
w/PjX0YwsH2m/naw+cG9I15lRRx699YsC143EVeu6PYQQPuEUSXwL25MUBvoTAMHsrQbJcvI0ttc
2wjcCyECsti/ccUXtj3tAC6V659heNeoB5Lk1AagOlmwPsd2DZs3ExTnQuvSlfFysZQ6qf1KTErp
GDmzBlIoWcaJPIuOpSo67ywwU1w9I0J1rtPcPTpCcX50gJ3Z/WWD2nBoQp3uP2EaHd8YVCV2i/g/
Pbfb1a4OVyO1CZVUDCYaiBaNwmw3Pr6eZtLN1IKboOWd7D9NSOvsNzv0qOr5vaa0PoWRGOFJxjDg
JQNQzTP1Y3aW7VhVBs6joR5uHaBTZVatFPy/OnAy770Rfg4XwfW6AS/fixFoPxgU16oK3dGrXbvN
uCCbunjiSkDcUas94mZdAYm4Uyb1OePM+pZuKH7oksOqPEsrFo/T0VFRfBxXCByCQ2GtFWdXSFhv
DeP4mTOhrhdtKtjUz5z0Az8nDdftvNaLhfAdfzJi+1X5EuaW75GCtJZn43mLBtv0z45uA0hGOMmp
PGRLpXOdg8pHJUnGz0JjxrjK3VK2Af14sgMsGjlK5t36mG/9jwD139MByLGR7KZUBEF3G+/gYQMW
R61G4DxdS1tLe3UpOHAPqZ6iROms+N/+WqMu8/ZkkHHR8s/Y1uviGUEXzauuUb0lU2jUA3C3MCkL
7m+/aNOujv3OfZkyfRPNllzb7EWEiRxea0VDm8nfSz3Fi3J1KAE19lHiDXWwg8jWcok8NgKZLb19
lFQqaeOkvnuBMo8Pxsd0MrGSrIv53DW9D/L+ubBcOcXEgTU5fhb0cOJPt2iNxz/7VrEnCENScW1s
ikFZOpeDrI6TgR9oukd99xy7kdS68FrWzD6ilc1BHZC5fFhl7bLP192IWb7orj2StdQzp68e7aEw
RoNS1/LWMc/Ms3X5jj/RDTL4oa5ABMj0dB+DI5UKWCjtwQJqcSFWcKDuUUAWGdY+PvXKsPEZ1xZZ
a3G1nmYG1acrdgg+qfQCr9vpueCFVEyCtBJu/M18yaLdBujGEierJQxkmSqKmGdHxFGolR6d/uJ+
m+Cq4bd5vZSvQGPrB8bS+XfQyxd+lFch+n6VrjeZz5+M3j0GSZn8xEWzpXn3O77QIg7Cb2WKVMQv
pkIFUwmbrM57os65yOjNXFs/KlwMUNmOmDeCMlwtn4g1C3gCNsIMhPDbAG/s+xOVoFxUX6pgV+Zr
2QyCXoLXv1BVTbb+LhfFDQunclXaT52KNVrBpVLJxqcsnJgzoafGftbxtmVP4VNS9PA8YrqPxMvu
gOKHBbxctkIj6NTbrq1HHGLRmOXimUwdR0pYD2mbMUzuOuOVTtHcK9TS8cVt2ljro3gyLmim00/8
rnZ6GkadGnpQiRJSR8AYqp4J1S1Wq61hvdRjriO/vycaS7dKtssTeIznsQTYgNTG0Efvel+NOLE/
mlbxzJcGfqToM09topEOUHbqU+fX+emVMa0LOX7BdVUqtTsiu1pd6lmn3hBCjChO4zoxaAZu57Bi
rnLCG2Mo634y6Tvt6vpIDvlNc3oiRgRDQHJ3cxrg+IPy13Cy8qB37NftSfp0QG55UIyOGMl5zyWL
/kSvlfHIK25wViVB7ilMuPYV2Ck434OBnvxOMDbFi6OdBF4mZK2kOOpmuMOLSE/UR2IrIgH8Jqg0
ysJoL43ZVWxXDofOGAk8rS+u4hK3oNHILoEq39D6/zEE/qo9KVGTly9qMmwTnu8wP+nKr2nszBAx
PxLIY8LqAkBf7lFDUyG40lmmGme7Ev+dAcSKm5e6EfuZ3cemP64izaMNKioDVd5CCZV7ciW+jVjc
ei+P/w3PgrSjFDYQoecP6DlZK/jrePXe87ot6VNo4KwZWBPrnbqgDTX49iY4FqfbLIuMeNDvrbl7
3rsoEFCx13FCYhIyL2WywoSFF/6iHahnhiBHjfiPowHn+URFWEgtxtGnwHiu9hlg1h6FdNfRieZR
8fx30/jjX6avjjGGTgbOHlWFaFkcWb1NUZIIFXWjDk0CKHf+zqADJACHtzBsZyKRbGEYPCBQ1YLH
rcfXrL2gV6lOBOpso18SvjM2esrXprYtm44jHY6v74xEkg3SoslQPv8q39an0g4fUtd4Dl1vR1R+
jIRD4ky+gSWHoAcPnC6wP1JLkV60RTq0ohHisUPRxr/4m+pJ/OFnFxNc486ZqSAsEaVmPLu1NHOj
5WoHZd4nOSmWl7Gyj8RkuuZVFpGb5k+AjciA1W9AJMcu22sBFqdY0kULg4Y6PYyHEUD01a36XvNk
Rw6dHpQDVdxNdkRR7UcSh9rt+c5ipXOsGTkgza0mfAoCgPxTulrSiqUANe+6/VGhcD1D7rIyBWVa
xK5xvVzS9eWLFyqSii4eNPjwTQrD4oby7Agh2dBjL0gaAbcOVzdcz9E0zYeE4mXhh1ZAkYjstboU
pPTLEx25hlJxSskznOP4FlLTUeMmP1qtUY+3Z6ZBxMrd6CL4Dr9NYuU8LB46/PIVC7uSqEVJSRVV
ioWAmi4NVVsSq4cggdHrL2vweYIzlYDMYqHNNwAAb1qhlM6XheXIrdze+B07HpiPArxBe+tkDhlh
HQJqE9RnQWkFgHyZKgwxEfUelYZZO1M4sih1Ap6yx7qHeLmeCukkMqrjeQY/D49RkK4r1OLusHYQ
SaC/gK7FKyRIRlMnF7g4g2hhvBVixFbErGb4kZBeebW5oO+bughvU6Y4qC4JPizN8OPenu91lh8w
wFkun6jqjw+/dk7Eg5dlY3u88Z3MtlKDqKKTIHIayUGO4CFGaOmRElSHR2eeKqMUdZFduJzdiiqs
eei/pBfi5SFSSMTSc43sU7V0pqKZoMjaIFcxztX5bo1PC569kGAIAsuVIhvRSKjZlbzDU/YkT8Uf
axBz9WYxWThDhfD+lGOKxFjzfsrKoKQE8wQoF2GgTTATk6KF5FXWBx618rDyXA0ropNjG7wBYVWm
/+kaM4hN6OrmLv5p4L9/vG16lw4wsZs7K4yBqSSmSBhJZyXJvCkiVdDl17y9SSRa2cQFqGQbdbjh
6dSv2jlpaWVlkiHIFapsM070za7U9thjePouCyxnahzp+DLXb/xuXfig3YqLEmM+q83XwZO01SbJ
1EOLLsoCp7BWKBys0RsGBZB9UZyuXlDlh0w4fii7Ru4BD7qBVne2TNmksFmRPZ4MGikVAdY9e4hI
1+7bDFmeYXEr8fvFYO1K8r22Dpe55c8BfX//84eKbno7nx89RSgPebSZMdq/LdoRj6YJal8m2oJO
aybVvmxE6OIJtwtmBenfwhu2dy33TFRNovRNcbUzQjPzEy2TbBx3KSg/Z5leIY3zjPZ4Uerp8SJT
H6dSb71Ph6YfXQ1dqikq0B5x5UItMdOFsjy3G8QWeTn6nt1kTglL8jannbGeDhBDK7IcBlWDfT70
Rb0tmA5g+k7FsJZ+AiFR5T0dW1dWUxNKZPRZn5dCZyOKwtFKadV39diICYOqOussYcwrmuGCs0/7
vDrYim43W6KJdqRl1JovxC0aTUW0+48hjjRE45BrxNXP78aQkquZSqvHZsfesevbh9+GQHfE24/P
z/IClMvLYPAPVeZm8OgfmjbbVpejG1herEXG6jzy44ckwdvSKM10zRF00ER/crGXZLUWFsaItH9m
xImqm8aM8TH/CepO5oj23lqSvWOeE6h5ElRGBWHA1++vyc4SjBpt6wIO0bnHMscqqdoKMT74abtc
Ii4Y7iT+c4xeSUmwwWnQRhZHcsutRgUdMpucLQHlpILeaVEfvDwgPnH2zoda946oIz+54SdwxqEi
QAfQBmU5394YP1y4Syhc54sheLoo8fOSpz+W5RRiNHaCwgiquinDXR0VjKVHPUPegvsjHGBMjXiJ
g9i/CCI+952IIpiIDw/h7WONUiiGZN0A43qfM+WzqwLopadKR/TohAJFxAC1JUFeJFlOQhlxICQo
hvPtsPFHvnwRnpmGlb2xtiatS6EnPPmcyXg3Ix52WvFV3+F97+9K124eHSEfEi1j9ozTxOa1BYwf
wRyKSn87LDiLh2D8ZfP3ICWL4B5q7LuJBVps3dga3YlggVP+yw2swDnZ4/Ot8LQ7+Rlmr49XpALl
oSGmXSkcOk/A32bj/PPKVDUicwa+5a4Yp6MFqDVEn/ZWB0LhdExo8xvc1oEkgLD7TQ3D4u2bTpXt
8KD96O6WPA7ADX86fWdbd4j0tBzaCw19DCbHRalQrpdjMJSKLr7ik2h7FnNG6nEjkxCfhPa2VERP
+PX8/3W1htXl+lEtfPzApZnUPWgKpb0fGz+QmD+G8YBNc5TOXsL81O0xQXitxegoAZrwHIGcdgok
DdruZbU7Udt03HyUdN05Lu7VzaAWaLj+Cn+NJ5kLKZXJO2YfmqnKUwnkH0j0uwZWEsy3Hkzv0KCZ
ZHm5dPSTDvHFF5K2HHEXg0BIWV5B9S1o8AbaUi841k/Rpyzy3nU9f6Oszggy/5Nec9tRXSr1OSoT
QqC8wte74+2d3+nDkbrYaoVI0wZgIZxE8+of/ML1Uaa08tep7K8WH5LNS42PEJTwDS6IZKLo+Kx8
tSLXSO6js6qkrBxUg7FbjSik1A+V/6XuiAeE7M0BB9XUsgALcioqCWfiBN1ROe+/1v18umUByo/+
CEaqFt21wGoy8dxSmjBRFTJY6gA9QZzIuGM3iEqOo2FDis1kLldHXU7512vrudVufAv8pKI0Fq0K
v7v/tA88/YkqCpatqYp+1XpB5p8U+hU7bC0R+v7SYZwJQkKFrknoiYholmn3X/899gAgvtc6HKTE
FgYprAill3Gd81ti69mAsjOns2+sVZ/j/ettjv8DIyUeLwRhkU9A2STT/nVZxEkah0Rp/cMviA88
QNNoHTZwM0PcOFdi2eN9udccy34LjxHAIrkWxDzlSyK55kRYo6qi1hpLQVaf4to63cok0KGVLnaM
3mGgDZDEsEvD9SEtYbRUrmYtFY5+rVpBdBXMw2I3oYML1V3eKJaG4ULHtYHXc2qI7BIfcevpG+Jx
Y/RbmaCto9QtEeBDHGgJ8NQcDqKrqkvJZJMe3RuZwy9DAecneUss+DSzNzmyU667XlNXkAg07Npl
183mWIrZgVNi8r+isRDvM0yQYh42ZtcQgyOwaVCRcV89AWwuJp4GpfxHFTPhBv7XdKhCV07IqDH0
YaxrjNPC45Nrx78hzCVNWxkZzRNYkVjEt0+nFEjEocMao6tBLtudTFE3VviiOVQE2oWfJcdB5TI8
FJCM+g3leWs9+XcSdguIjQhr6w25y8g3GSCKbvWbNSue/Qnq9pkFFBL1WyiWImazGYf3rM+PLxeE
wIhIpVPAklnHmjaYKMyaMzJOND2gWStP81U6KzelFRKM/+NOn8KHz8I3Ghzs7mSR54PE5iFGvFkN
7tYN1PwcDRUaG3Y5AItJixfwR+s6rsmQDSBHEsagQZHxynwrdl9FhTBH55L0T7vIn57xGnUnOXyc
S+rvzlRKRDcrCiPN8pSUBFdSeeTrgkFYspUbJmHNeGmaJCbXA6rtJ+ymUPOV6cnWizPkZCR/hFZm
n76qjQmJ4crBGspdpwIW3gCYf8rP+WsW0iDNHTB7bK4ytBnoZEnqmnAMmOpMDRmVS5JKVor9UmUT
xoweo5ptZ/5V5VtMy/LtGs7jK2VuEHgskdCBnrWWDB0p23i8ZhzMx+uBT9SB/31a6EAYgZTuadL7
C4w3Mx5TpqZFObDVFqnIqZZDc9F/nCQYGyNASjtojm49RbchFmPT3DiWo9S1w3lhIGHA6fdFMSqL
P9fsYeaGPPjKkBf/j/UrQmn8SS3D5jg2irufKVHX2hpJ6sUOhJTH9JaizOpz/LpmhIGdiQsiB36o
No6s2rGETlonmkPCNtRtNcKJCSI5t4kKTCLJwvrlffqNM1GsOygkNQArCvsc3d0MJoiAohgLr4Mn
gqfZYwUvMak3eVw8UiaCeKrh6kKm3+1MPg0QekHlg/FNN5rnKOvDUhEKVqMECH0VVaPSwYiJDB2O
oUY6xH3VptoPUub9rT/Vxm5J6BwXH2vKHK7xOQC4/CeD5OWe7QUu2wzcWGpwsRyZQzGxHBV0srGT
6ffZsrUF70QA0TAzJ+PZiHE/JECcTXQPGBfpMg8lvDFy7iIu4Yw/usuwNlOKXfZyGvUunZ+SgJOr
cecvTVyBvWZ2Y6ednznK9/utsd+zi7A7cxUV4mm0WwqzX/RUx/OrABvcsbqlbrusRUEpYtBsBr3d
oIE9j49TmGwuZbzCBKLGJVgivR+3YFpv89aqf3o5QhBMhLAwjE4IuO6yCZ6NVOCyfvIOpOtWAMRf
SelpLB2LpmdxH3JaAAoBPEiRGcIv2DSWyBdIFBSvLrgao4o5fOclircl9YxHxomalQK6nRaSi9V/
w6Ro0MD/N2j6jcwlyEdfHjRdg38PmhGC3+oGzOszhhAEtz5ZphzS0mRUewJeg5dV6LakqOKA28OD
2N0BKmBUw3XzZo2SWYw7R/WDGq5IqKgVebxu//25niImRFd/1X/3wudUoyS0r55A3sfl+jJ6Vqjq
/1Oa3tWXYdS19bsnzgy8AW/cCcKPUVIuQAraMZ26YpUChLz5Q1wTywAeteyxFXm1viuuhnWuj2/w
3KWbuvOvSbijWhY3MIXqzi4IAJAqDtXe1nu0WXeKc5hnrJ2ntQRcm38nfxapC1grLrO92iE9Qu/r
l56vWZyJOSM9spk+YuOuu2VDeXi2VDss/6g1e+6iIZR4kTXJ5I2vHzPV+L3vn7msKDpxeBie6RQ+
D2SZqdKnE3FaoXRTgunoIqYY7QPXUgW2S+zI3AYqXK0OoyV8PfX2FoWTRZtCJ/H+t+12ymp2TH/H
KlYkffBU4lcn89ckKj26HrzL/mx8MXEyKzeSv/3Y/sUjsemqKHl9Wic8xsvzLDEXnwaXlBpK4eXX
OPICYuDOUdIHnxgT4PYTyL6VMorqjPNo+90UtWL6G494qPqO02Da5sDM7DWv/3yJGEdaDs+WBPr8
8N5AEgJQ0gbTSyTjwBdDOVDlO8iqugkSg35g7v71A84A2KJ7CcDeSrVPylRu0d0d0Yw09maHCi5I
lAjjLlL36S5Axt2Ey5YxvufYCLLSFBNJqOi5uBa6AMfQMkYJZt+B/wslATI/0IYKX6KRIu5YPkqI
MzyF73HMvFaEc6YsDl7J1Fd1M+X/BgkxbI4DyMPyaEFHIz0VQoBG0H2mLABKASHOIQIfFWeRkp70
F74xm7Q8apg4NPlWfEX5JS7cDfg5uGBLGWwnR8uwA9Y7XPbVLOEsbZSC6rquXOMw8/45R2M3oHGa
f0m2wEQtsgY+vHIVGY1BcCwGU5IvIwB1jRw+4qhc9+F78geG2A/RRMSL9+Agp0nkqCZ37vYgzDSA
kmeMlcWqhPogeTvCarOA0VKjDBXMykrt+SMOb51mOPRRja+/10x0+QZYiusAhvb5w+SJ52BMagtI
bpduVB38sHg2fN9c3CRwBZPDlbjmv5WQGY0HiJy/EkuHWC9Gj1IBHAfBGfkRKe5jk6nyoAyx3KgI
sDEROndHyYUwKU1s1fXE4dyrF4vD4G8ZNWR+HARQ4+Xd1pCoDjuS4LYl+UOwrjVJbTLyydbkWazZ
TW+OQc+s8+ugERa+gV8Ne8oNo6gzQ9l9SXf0VyiG53HrVh/EtYyKctAfgikS3RBp4kc+C31t6P2P
wbqNSbmAa278Iiyz922Kb2A/lGzbGAodjz2+KTIJVG5tYLFHbX8CkeG5rdbXxqA/vsKptt35x+t2
5qyILNRHlx1cR8dLQlHV5Kcf6Rd597Bj+4Xwzxhlg+HbywLyaWEk/DuLtzpKopOJw1QLF1k5FUxO
BJ7yJDE4ok3EnWVJQl6Ou5EpqMbocJyIGO/aao/Vr3OXgYV+U8u7dIxVm9+5KHLEuwdUFphmypR0
CjaP3DUTz3SXBofr33UT6soRpZXM1mr4ZBhvgmp5A61YB1WkqgYcPW+UNm6O6FN1WJ9d9juVnH8T
rDAqCJwY1eC6OnopPXvkQtHSVkw72a/BFNDH02zl0EdYYOPFRD1YjOnfW6SuW8nn7Ff/uAjMr/Zq
QYVYmTjoIuzPEK5agA5H1r2xM5SGIP6z+VtluYXyqJqndbGgmJ46BrYfyYSzmlV8dLmzi2On5SPW
SR1lIaj0IVLw5D2g6urbI3KeJx5psV17gmtk0pr8uACfi+cntjUdVN7mRLO1RoGAExyIOsVs1Avi
sx0LVk5BG7yuX1X/2zta5tQ14O4q1QlCSQJtjR9ZpUm4fxY5Gia3koMhtL6pBoYzjYhRtlVvsudp
ldgFBmuQb7GmBHtLvUOl66euO/hZmeYyCuSV/pWRJSBzUC8kzAjrHXI+Ke3KykBo+FkNS3Kml+yq
4w07KgjfMgntVn8j8wuWueK84kW/Sd/ON40IAW5aN6Mf0xhXzzaZ/Bi1QVr8F8Oiw5hI76mhUf+/
tDSldf8den1IN6ZT9C19F0dkL8opph9o3elgJVNumrWkUSBMsFWaRBtPe47J91KITnbxWP87Sedb
ea+QOKJvwbF6xSNaWcGnsSR13rNoeqkN6bOLMNqzj8YcUcMNHoOOxO1M29qK78htMYPhy22hFiVI
nElfkGzFaWE3D/ouJjDWfs6X7L2Ueb00mrc9QkJIrkO5boI6d6cJx4w9XxY/WkT+iAuM3vUSgQAd
yBOKOifR9bFvpxCEuyRLwx8dKSWTxLNWdLWEu4CrBJoBcwQQNxcsxLRAlV5whLTZUdxh1aNqbaQy
tb+ODRqbZWazhR/UOjaNKnPvwgLiJCUDGDnuA9RXWl6IfVUwJ27syuhCgSmNMVNve/Iy2zQ3Zc49
HD75Eqjet1kgsykRzhFKO3LlBLJ1OHhbcdlNFS070sZXeRY9FOAJC3tk84Y9m61+ZwTlexH+YqAY
BlSKKwaijNIZH/PqorQVngINbyXMKWYxNav00t1/OtpOqW47nZfkfrGrLv72+PNyDeTlBZAXJpo2
N1qeL4U2HQ/PVSr0zS6AuAfvaPVEO4MCacUTW83I00LqLsNcZeDusJ6zaK2XgEHWO/E5OS/ysCyO
6S81tn1KLWVkUpHjTrYLHQ4ivbizXn/zVfQaB5P0S6/U0fUzDa8rwZz/2//CTRjpavEmmr5CEN3+
kXj9fETjchcxX2ODyIbD0aaiwAtfzAQCfHJ0gnojLSMl52hHFTbAgUgl4VXpHYnRqJVyW166jHdM
0ESWFWJwkNAlo3VSk9Xs7v0R3IRCyN/S8+o/0etsUFxrUNNv9p+FjHqWJM6i2i+ZwndmcsAlHMrb
BHKIKGDEpdz5jX5Qh32IEcaVYMUTvvqoFjQqoBn7TZBNhNARl067LLU5Pu/TJJ/Q4m/wIXW466C3
eNgjLuMe3+GgX6A8fwImJBOEkjkqpkSGpaklZUl4bX0x5E/33jfLLqJMt6xrESpfWz7MKJfpfarD
NjELcfVbxIZVHKmA+F7W3uqji3MqtDqQqb3O7gUWrHFCl9oiL56R2zAHxQ4/UzSpJwUfd7Vmx2Ub
gT/QVC4Gfx8qrXfRLr8E39hyMGiqUgJYXZbNOdge1lUeeec+z/khm+pf6NZ/g+Zf5ao7Ir1AYyCH
C2XHiD3NX67yri594LyXxwDHqHTE7k7vp5CbLFJRjDOhgdlIzOgLI8bi/6iuABaEs9e1dCX9kj8S
5jXJ2CyEkG/zE649KXcuIuPmphj8Rkbled6J3EHa6oPSRq7toXfOjjHQ4+1reKAPuhpDoWVkJsQC
w6N6W+9Kv1MHskldaRuZ2ElFLDWMYLjOjplJy2b3qzcZdxHgP064kbNSF7Uq4dE7GvjA6lRx5Nmv
D72m/Bpx8W2xhk3FSisiQ0uYUfLQ4RoFzqGHxEo4hn6plXlr3gxCrRolkoVR2yuqWZp/e1LlxNsP
Mal1we+07y/oANmRWD5TuscikYA/scZ34s5YSCHQU0fPAflpV90sxeVMxq8v9ByzqFyRrFBI9sFm
FyyypbVRyoChd6ruEeQfRjE51L2fRFZuQfAeHoMaxwWSRAusr39DxiTgEmH24TqsSfSOiY6GQp1P
LoN3RQEQ6oKep71bTMQ6NaVlb0rw8EMPOAPuS+fuKLQ6belO5hSFoOSXGTOCPRvDx+XkWHVd4kc9
Yv7UsmTgKXzLW8T+/H+wShl3POF/bUearHT/xa2jPSL7glPGUGf6RcnymghSFNol5aVBtxp/Lu1S
I03yhMqMyFjwaPmPEhe9M8CxspRWULDfaCyRZAABxEX4f+BCOgGc6LxIbE1JnXcSFb0LfTrFQFnC
ZNxCnge9JWcq71XwLbQ3F1imYWMuQkdgIkeHrvzJb8RI5U6ckOtvn1JZArQDnjZ4n8vrrsdR9MPg
xpMGIhwzi8KXN7hCLRBRvenFwEWrALHxEGEDsd9yIc1kZVoLeT69Ceow9KxdWPlLEdgjBAqLFB1c
zBpoz2CLfTcgbi7hy8aYerQ2EDg14f9/xm/4cQccNnzMIhhthqrx7VoNJ53Y1JH1TB5RJo0hs/vO
cPTjHiI5mH67zE32+tU5EtoTb9lr1zdIGX/v0d9W0JqIBWx+I4lQMenXTVmvVkQT8Sp00nq8DxF6
F1BiSxyep4hNmhCp5xcnQQ8H2QhIvTVysYN1CyZ5xeJhOBiSrK2WsjCeWUzh3uca/TTh6t8wjllb
eP9e5+2mo5X3/rGwBzSREzu21FzQ6JdRSOXQLvl4SDdQcp19Qca0wTDTU7pfR+ITJ6R6rrH2hBHk
AueFCgsfPO5+c/IZjDwswKocuFzCiyXevxzaJDvjIlqPB5pA7o2EMbiY/jxlRfrFSJdUqu7KLZSS
weNyLaejzzE7tuqfawql5hsiUQnKBeW7u79CKksC1poIwma5k1qbxdcwMvqxFL+zbdm8sNjgovC5
VQ3xD0CZmxz4rsRlnfQ4c4XpIL5fNm1Ki5dzTqLaUGv0CIMu35MYcBQoQh31jvbVh8od4AtoIcZd
FuYOD8bQy0VAJ1T2bYqDCAbapLYbET7n1m6GooZhAm0q70Q9MQTwQqx3kLAu8rlCogMOb1fVmJ0Y
iQ4tsQFLyKPTVN0GfYCPjdrsk43RsLEeF3h0YLtoOuPQ51mDpIBVONw7oYeeR9owbbqbQOXy0rM8
QBt+Do8vya04ySB9PQoCqJRCkaz3zbmv2l8mU3NlpV4yRcjT0keC+dx4x4kCg+eq4Lx0PM+5O/Br
olfMB+/GkUrT9cXKWP96K7oqmlpWyArMdW7lwhBKOHhrx5JA2sWpDWRJk9MZkVs08bm7NBMfcRwT
PBYyI4BMeyix1ZX1dFreqAX0deONQVXx29MTonT+ZnZWbNtlMZdPmd5WMZIzvX06lM6U64n+rixd
wTEGVxtD3scqNuOXdPpf9gfJTpMxKrsrBdfngcuFnewmsYqV4shnpRljZ6XzeWU+0qxDBMDoXvy6
PvLHPdwHOQGGGQ4jz8bh0I/eIERU78CNEX7Ht1OG5+8FjZqkpYAN3E/MzBh6f0OtNHbVLLsTao7L
zkLHDH9K+Uksc9GGVUNAFdCFg8zmflDYySXDOSJ3AYeESGZzfofygBfLAW2dYun2JQPn2UyZYbIw
Y/n0T5FY9tl/TAMBwPbeSxWjIPY+AJeq2L188AGASN6eRUYIwl78OLyJZHzGe2I+NUorXW2FEroG
uhkqM3nUF253KknW6MNlFGX6t//l2YDvDAgw9/w1XeGMazUTUV0mAdLgS0m/AR3oOqeLWgsfnXtU
FnS4Y+ZiIHwubnqxQYnbMiUX+M8F7r8vNzjOOwsAkZbPSDSCBCM+iq8pcFJj4LosT0RtpSeXak8T
/kEObQvpGcEcIt691AQq2nFQhKylkArNN3i5KbiL78wZMjHC0roEnSAsg3m/8cJT/rDAo/WczZkc
E2SB3KgYn+bMEbjy+pfTDU+zZgqPlwYM59/ryMKFURW0knucPtLT6NUx6rZ5lsxl4VcwRKPCssyo
Gnbsz/j0exFeZfmSr1l+IJ8j5q9A5+CT3GAJkDPJ4m0Cq21VScLn5j3cYw+IcjViSSd596xsFAje
4ygsCEQjaikbZpM6fl18VMnV4gLjnWkZu7jc/wDIbgxnRJz8ndISKYfFD0FaRlZaQQt8YRyjv55L
ZpLckvMvpJjAn1xk1DC1A3Ksy2s5z3MWJSvVOIRlm1iOcucUOCwKKwlyZsBYnqDGYCJg3WE3AlGT
mYcyZyeoV2xSgDSoIXo6vhIkJSwV/ROA6K0pHNHZmRL+AUNwFl4xVPeM/uEiu21/cfv8IgcqNZLB
1NLF9iESWBrm8h1DQtSzTOVJ86kzN/Ckv3ZyxaelL2r9rLtmdc+9/OF4DpFCbnp1wjOUzufzcLol
tCics8KdE/gtYQ8m+Y8SN/Ec5IXcHuCyJiQj/SRWl85JPeyrO+4jtnwSo7dEqAI3pUlSN1l+k+O8
E3js7h1r3xCbkCZKZDravMJmjLp01qq7zbFmpn+gPF1NUtvJcRO1pcH2FmkF8js3jiMnz+jzB5wy
cgeFBiLiToA0GP4W0xybxvL4yjAK+nvAtrO+nUjZIwy6HwXLtt/MupDrJMncuUD0bknLpWxXu33L
IZy1O85OAeFDkkJLOuvFdDSQWILbzCqLatFOGIkQiIBZc93G2hUHTM7q9ntxl2A4B1g/G2u1A17+
yk6vmiPnHpexTL8+QAgrxU6A1hVcjn+2LrI5In+JHQgmGFIEqT7fZam8MKJ0k044z6iaNO48CyWK
7XuXQ8Gz1vgzUEqzYb1bZFN0Q0bIegNPLIyq3SfGCLkAutZGldwGmApPPnPWk19JX8Kjcy9dbQwO
bckEvTAN9ZlLHIFby5Bi31gzapIyBwjaCLcpZXhHtFJoTWo2C6QJltLELKG2EGeJc8DqpmJk2k5G
iTKlS7Dl6qm/5rbPFrPwg1jvH1tkq7rPCNlqL33jbMqAczBIwq/G75vBFz95wszCffp7bErQIl+U
w2YLQYQleVPix+v+/qHtYc1D9FYkQmaJtJxbZcRZdp1KkRi9IXyhMlrFBMYOpP/+FQaGQMoBddmL
jedArWm6iPG5YkmvqQoB84o4QlVp8IttOf1yNS5Jt+v7VYIlph1Vev2H+Px7tj2dkCArWIzUb9hJ
3I0Uy0i88vgxplht0rvCdaqSl0utoTGr943FXtQJr93SaRL9vNGglgxQEmxZC7OFpJkV3WlJw8jF
IEBEZmL6YuFIOijtOWErJviiKRdENpQI7FA9Cy971z9jLRPrBxNzLmWIMyG+BaDR3WNSBb2F3gr7
yuZi2uC7qSKwYhiksKcgwCZ0oT08CJotKOoErZ6YiNRFyeGWLVwbL75XjRUM/1zo/Z91P73Qxf/p
NUIBy2MPMNi+SN9VcwTYfU9Z0DFcqmzSzFyEAy4wv3a/Y9IGYyk+uXemYx0winm7NVxiWqYwhsA3
zsngcHNT4sMoO1O+/sQ1ukbbyxjX/qyjspW/ubiCsjickrkZxFNmKx3hKr3sT06GJGa4ne0QAyUi
c5G/tHOr9u0afPiM3alFGxuP6cPv36poBJOAGVJYZCKvLRbmRzZQlndb3lyOrpwJF/mt1+qmfQHu
5FDrrLwcbgnHxddtVj2olUCgelb0CR48uD/MHYu5jHliFdVXe6m5ockBpVdu6voJh9AQw+tWD6Fz
zYa27qLVo3Fzf3+Z9gI13Cu+/Pfy4BJi3YovVEl/BIfCXsk0Fc3xCgkxdkWdA4W93khs30z10wc4
w0M0W+/nn6Eg/mpaQhYj6VV6Ahz+euDQUKojuBP9LH1pl9kfKj04VhQRYJ5MJ/i9EsQ0jD4rlOfT
PzhUWyz4aTaB8mT26RQRSzrxkRWByQG0XijpK26yZRs+39URPtmUP8azgJHAqjjYR/qkAydD+6rB
eYJ6cDnvpP9hs2KcQ4urUdEyV7vimxSgYyZ2R6KBfUOYuT00nE0UEVnMZAwpWdKN+9fGXTimcIsd
JsoEl5uOpuLU89xEr2Xl3VlBFy5qunYZVTF1BDO2SjfysoMy/MuAAVa4R9AUWc9baBMdqY2mlSN/
kPtZE4xe82z5G9uuKZmfVHw0BaSjUF8t5jfFAWZf8EvSYqc4xb9ROlopq2Zn5iW6kPzGNbYU4C6t
tAKFKlNhEZZ0oxD7q5zkGYJHjNWVIT6WmOUhBzlskmqx75WLxBrAM2DOisWarFAi24R23MXqawlI
Ai8ZUWqQbRRU8uqR7wnfitkHNKiCuKtVlFz1HBbt5KvjR4GrzCqko4JIErvmm7dcHybxvkyhC9kr
tk1IpxDLTtzObvakwM/o749rU5Y1bxQb03Wh9T6raJGy7U87K8d9a3upOBnBc23D5goH3Id4j/yZ
Jh0f0q0KdyOYtV3jc35PWeaqluRXmPRTHyp/pi/nQHyEXkWechVgzyWfSY1rprkjAkglA/AWTPey
lOV27giznzAZDsBAkOXN8zugrXedMJJamjAhVL4V1jvNkkl1RxbOzUNFCyXk3D4JOJ4HYuLc6QVd
wcq24ffffoKkPgmPrAe4SB3U0MA4F+3IgiU7kuLaNquu1AHi0hxH5mJ9LSvV4ZtDNbqB0QfzoaH8
CRTdzbG6ffJ8ctyNr/NgWz+6bUHGL7P5fDt8cOBw3XJra7fxggRLWpYaVRqkEiq7oimCWBrIicZU
84I261kgOIcpqGP7/nMKPNGva/5XhWl2QEXmtAns2vAtHNB08siynlj4DyKpoe+STnBAssgzo5mg
sv5YA55BVat10Vp5WnvvjCeUr9RHIuiiFrfz5RAqb5E47B6DqE+mQTudsaMatoBq9RFEwy6u6nIt
xE6CmeufIy2xheuqojXHPHD0k+wp5+gaJ4Jm/he+A9bTyNa7OvooNY1dNGF08A1/x72yTmf5uzQl
3YF84AC1ELFIe0WrdOqspQ67KqirMZqmd6h5al6VZDmMe2E1UeZyR5lIXToCi6FZsGIf0OIctMGY
SmS3NzYthtt5Md3eJPfGGi9QMotfNrVinvEEFCiuy8GzuMRP+JRn2OquDrF3Wgi/jC5/WxtKt5LW
UX8hT83LIaG3wnh+5C6XZuLio/1T/79OOKGoKGXMYQsUjTVKvL8eSY+HGXZrBWeSuxChTG7L3yMQ
xIrFU3uGNGzRYQTbrLmatZ/w5sUfmbzijxC+8EIihaJ4jiTJ9xCnv/CfPDD/KxmaCOOy6zvY+WyA
Gk+ejlpiXltnsWEMpbKEKz4GwVL/xs52Yjk2XcqXL5bUxr9c0khjkmZLOlwh12TprR8imhaWZXRu
GMTcvLYpaEZ8hgkQR22Y8u0UymyP0Koq+RFsOmHJntUkHAsxbwhm4PeA0MNsd7mSuHQHfJ8L/CdG
sCSRiPzE7x3Yoo9NHevGCz+PQvY3la8QdAG0qBUxIyJCL2NG+R0o1WcJ/s5zEa6ax/d/QNJwuuj4
hjJGjLEYW9dX3V0lSHIu1mppFxKkgAMDEBsSU14xknJLZ0t2h5nLHRPeYsw4qwnefloiFd4WG1xV
cbo6Aj3dg8SCWsT458+I5xGfU8NnpXJz9OLR74kuNMYt/3zrPTPeyUpjsQWM59hBiFRUKFwY0gB8
Bbezhjw5vg09uOO9PtaFCodua59vxvGLbZRXy0kIJ1AY/Uxm4tsg/Bw1PTo8wXXnozoFkR4iboPQ
xsiExwD80SJEDNepHxyNpbMlOi4JySzm+x4jKz9bErz3QJE3VaeDoWxyahxCfJslSAis+thghwrs
BTzuNpIwu77g4XFmBTl05D6FISILexMIuNN77ALsYbD2Ryooax/iLGIrEBpr5KMHNSOBZNSLZU9t
vI+uH2KROYlrBOF+PFZDGCqD4GGkmCsVH87twnn02LWlQXoJ5LnB7kXoypio0D1v9YqjCunQJSBt
HL79tKBPS0ne3mFHSXC/twrdvecBAzumPi0cDIVMz7CCvF26jkcoyB7E1sCze4M54wm3Rx+PNCMM
OsWmKTbn7tbL3LG1qfx+dzGXi49T+rLM0zNTtgXSmj/tHXOUa9bBmRulg5JyyfIgvjYHIPiItc+k
TLv981wIIRJS2PNtw2S7ExFUCvhc8Wq/EGh9gih9UaQRmocibmiOjWES7wJF5G2WGwnRMQeyqxJd
6fJZoBgu90nSz65DlCE+iIpqsrGme1W0EGhcHVxg6S8eUTj+nVohHCgEzaefkw4JNLk0xlFHm+f/
3dxCpcG5AIMXtWsjl+JYh0wpGhDeHaXnv5OT0KArIpAji1o1hd1L0Ld7UocsrNLBbMNIyRlqqBxo
Lr84X0vERvKTv21Dl5evtasHuJqzwlc8i2OZ/lgXmPjkaasS8aMn8YhSVKKiZG1aLT86LrvShZ9m
eZbk1L3f2rfiNiXn/D7cam3azrHhv35OFmODd9qTahyaZ2mvrKCbkdvZb+NMSKa2bF1Azs7tAbsn
hbCko4I9FujFm+KeVxBz7oG+tp7ptHHCCTZ6OKcV1YbQjwafpxDQtw/DE1xQPmeDda0dM0NMCKZc
tW+H6oW5VrlZUgHNaUJtFgyKnd0lRQPvfGEaplVWrCX+MmMUcJlP9KiPohFVszzyVoGFDzut+yob
0bK9ONk3wGng8O2XVz14Wvi23ewitsKY2cLW6gnvw0PlorXRMf0jNX1tWivzvQin1OWA+o7KXkGs
cgyywq9z776o43DXQjeVf+CUbHqw+JTu+2eoabwGBfnirniRQhSV3bQuXUjyHTjAuVnIbNWlwpsl
u6mICpdy/XoqIwOspzJjrA4efdET9xiRWUWTAur+BWpR/Xe1YcZRau6BfyXG9V6D5zaTeJURHPgG
8DozbQ2G3odh6skAqGvqMglwUtujDSIKPNozR1T7NUe8Mv0HNVYniiTp7fMhXclmI3v8rtvA0L82
4+DaJMIZiWSbDa0fmQTxotq3UjY9gNcBw3NcAPGL4hAwwCYU9gu/VruckonwUpG4u1gGziEIUp9s
JlqZ417p3mK1riU1+TEmfETCdve2w/OhwLJgfVGnx3V6goy1xnEKms5QSPNefGV030K9A57Nh48n
mTzrZtslLCc/a83Pae/4IIuyLgAjy7QT5i11zLFJgdQG4wf4BRfi5FRX2mRRZYjqotan4w49JRlx
6XXtpr1MfhYT6FHqop/HdVpBjMJRYalgTRUQ2GpluemIc/Qb7rG2afW/pIWZDtnRlPvgpsYevf7E
bV95RyT/aAr9oZPuvcu30flefhgV9ikX3uG4JmXmmMhs31n6cNjlNaf9yY13t9FHBTG6E6x4ulay
qCqYc3mDF43hKflqkyjhjD68oGddV9zgGsexvR4ad+wCQ9NnR8Jmmysi4twt3u2XjiFkgivDdVG4
DQw09Y+LAxNyZW4CoBV7Ou87mbTP5Npt2P44/qOJ7UrsXF7xyyREcTJ5vvkoxqiu0tESOt3pG1NA
okzCHJrr/kQWFIAXcZm8ziJV94i+GMY7bJJjLsrSAlWbbt+oNAhSXo4QH4ANxbrhtKwGj1HJfykf
6ZrhwyMfayj9bCuydOWhg5+hOxC458sBkGvX+0f6kx2OqASs5+bXND3CO/KaIq2L1bnSJsdr2CIt
2CuAXUOQv+S950bvwahrWfvZeKOrdQlgCtG96vkIhd7rcNE5SWPIWgDbijYY8zncE3Pta6GkQICU
oOQMGGr6hYYuxjitALq5gSPi/j6YxLsY1P6BXCJOqRH03u7zY6agIjh0JGS97mQCEFVBcOzsQA6I
AUXMUKgEkDLGhwnkAeeBb1gSqTkeYp+n1XaUy/J2RJGqFoZZY2y2JHk+YS8oAr/wknxHxYrxkUlE
pvIfzic+ZreLBFFtrvCR1nI4iZR66iZmgS8UO5L9fCVpxjsi60Vamh0Nz0dLNzUIk3byQGoRXM/P
WyvmutisIXMZsHpHMh4lWcuQPeLBTc8uiRGnkCwh77w1TVATVW9yhccgfp70q566GC/zjH54BUuH
8BGA0U37mwR7QCviIx3GHWiezhEvg7L6iRfIzs1ktvw9ugLjttulwGs79jQHcKddeJ+CHz5f1Zb0
T/sfL3U32LWVRxx5WJh+3nrgCnPRjtMzR7WipJN2d+Co49mSECQ3H/tiiSDTvwgJN3/q8BheunL8
5GCh5X1yt8pSpdM3cSD6OL/drtCnk6hOCj1S7nzfZmpjZP3nm3JDKm7SqEbXGLYl0pGfAIrFfNkl
Nd2oTqMp4PMJdkbi/jfQzQOdabYTBqDlUexeQBcUUUgCSGPPuelH/CkO+VB0uD/zBPkNXiONZxhE
iBpTIi0l1YuAAt/CdhiVJtIzMdcn+CC6NQAkLFhVzodsObjlCVrVDjL5QY0OHC43LwMSkb6Smn39
tJznFBrmJEuKsvvM6oNnmoWSRrzgbtMiTjNSBrpC2ChJ9yztlhpLuim6rbOGCd25gMN626H0UMHb
I0kg2UUlfTVyCifsgIR0/1WBX6t2eQzTYIKUagvthALOVKO0/3Qg1iNas/d2Tl8Z79Pjgy3H4O3H
ijXQ65IAkIfKLZXJJFzJsJlYYiDLwzH6A/kSJf76X7CkXWxsIhweKgbI0g9pWMGtzYSj5AmFV3ZN
cDJvXNXOiakPAKWEQ7DPf+k5wpqWN1b3Klg3Vj8DcUmM5OzePgPGmuwhfMuqhdTv9Xx/n9CvdCO3
A0iws+i2D8nqiwWaTQqlJZ0+fMlW722xlBVS0Uwmv5n10jJCaye8ihWbhdHVpnlB9wXReIG+qViU
hpw3HkLtG+NVUGUo0/gqigKY1sxcmTn3OE9B45FiO16pURhqhnPexZo8X8ldnrBFWXE/BDrb2HRi
osyOxMSuR7he4yQjJpxd8Bu/Knb1/uGItnc9R1vxCA2WIM5yfM1aCM7eDI49t+pdRuUSwGy1qzcc
KhJoT6CEwTDZjILGTaxjTA6ncIk0fgI5EB+OeDB7cpW+QHZbF8L0dvzbdClfcjOMsx3ofFLrue7g
6BdogBTpt1uW8OW1HR3F9sDT/NjMJMBpiaZm54nhYyHqeemYyGA1BWMi8eBBs4K+Ufpf6fORPC0A
BtsbAEWUIXi/cq/1bpGNgWSbTg8FrNrM93LBW0FGovg6Q9cuHj1HLvMuihQYtgbAC/kMPUcggXkk
LIbNpo3kBCk8tA4/GAoZwsB7tHUgQy74ajDZSBsvMeySuk0qWDPsiaDAuc1fIf++Thk4xF5KD1oT
guPvPPs1oEZMiMaaXxlXT49xdehd9zp9khW7mtIMkC6PQil2I4tiwyz0yABEn0KvqGpIyQ57nquL
mcXz077ge2WGfDY748PkfGSxFEiIAVIyEAv/1ggLiGdqKbg4/kdC9YgX31xVtYZYkhGgl7DUdDQx
ZArkpPiFGvTflBG52hK/BsPe1LNqDl+OZrjrl2zCLU1DJoDZ893JHY6/UK1hdP4YkdewFxg3dCX6
9FDSHcaep1q+DpLRS46HMk2v/ZMAtafwOgZaGklveBeYS8rkgvrGKokC5ecKqQqAj7HBAx5hfC7b
1RMcBeEtT6n/4h6VxHo8tU5sVIMuV7eu9Jqp7/Z9knZeDz7HvL/5mwPN9RA1DMwhbPd70HIaTHgp
+bz/QrXL8wJrVv8/DhgTibAku3nmOgQ15TlsCRR+zYUVFTWWrZhuwDDYLbn9hrXPTC4qvtlpjTol
bOy/2IFEryYxqsBFHJWj761CioCZFzatfqe135vd7dxvZJ0YNZ0ttYoBiBXdpwx0CKUOcTHRUsWj
J4KUr9T9Hzmik5YBwb9KU4RTV+rhaiJ7q2+NOj6iu9+DOneECYXBRUVgsLGr60uVfqm1wkLyCgyG
C73J0uaVxrr0CKuSlWK1FWL9iiWsarkiUwML+gz6Vrt0odzSYqMwwvEpgjqwoh08rwhPpMi9JeDW
et15PY5hUit9wYQ1Kva43Cl6BznczHDOdYWBaJw8c2EjqPRKi/PC8OsN+0svuxUVmtbRsf1IEqQG
Q+u5llcuGfYOshI0VtxTf9Yho77yMMNHZXa7dnHWJilzs56lquYHAaXQnTkcqXxy8c81oDYaYm7t
5Da1etAK+uN2/UDxWbgQQP9QG+EvbgikQSzTsSSXuHEzXE0RCVq1j16NONvVhw4Zlmm4q3cedJ7X
N/5BAhrE2jT8ptDaA5FHIWdodgEAzCjCr7tbcJhbJ+mX1t5K1yZ9temyYFKTAiAIxdqmowD0E8Gr
6jk6Zxvq11APPvhLWMSY64tdGV2LWe/CXSP4hxWpk9YlBXggWJdP+gxZluUrXDj7XmfRiwJAlIUQ
TSt6+nWCSmrSDKY+e92SY+RcPvMcdSnkxm+U4TJwtsN8Kx3CuRTxmanuBeeKAX5SBxMnzWROX41O
u/VGFHMUug+PbgVw0W7sf+e6OMbwSEcevHo+uI5I4POfBTyUpdL8zqkItpFY8sL5gIQmkmAgm6kI
wrwkf6anqomJegkN+DKG+FlZCVKI5h8PqkgfUGS2Lbbw7rEnTi2rB8Rz5z/Vip7p8BPbeBg6Cfo3
+rKQh4uOP8ZzJ+crwwotNQC7y8cxMOyZfpowI1V1tYmSz0mOwLeAuVeBeffJuzywNgB8+5AXVUBR
s5s+nOhhyeLQKRIo7OSwrdEtFYd20w2IUQfXvtRKtKxCMfnJRNOS9xI2YHTe/C23YsSQuOqyG8TM
M9Jl4eMO2Jkleu9FkXnPA/Uz91QIvGHcRafkC2AoZWkBXVSCANlzR4Lqq4DMNcg62/Nb5qq1cbMp
VUYw7R46GA7aBxOy8CJfnbuuDVuuTu/QHvtIYtyQvJCL2AOn/eSpn9zOSKdKnq9qLpblV8jA3Se6
saso/9BWbqMDEluncr3zCDc/UUTfUxOI3YzyOTIUV5Ps9ede3+gXk2Zhc0PLW0a4dsNsOuQ/qAzF
IhbdMz1lnd8hGg+9k9JxTNJODGEpnUN0uXoDjziFwEniNMOpqfUM7or0HpTIf5NqNcRDfLzHApLC
wMewAQzxp/FJ3mBOaW3jDd9Hy17KBrfJDY2iOQ0rEPaOH4MQNz7WlYj8A1eiYnhmGLYkBFpnY0UE
0WwWhzqMLgniEP5ozO7vuZ68QvUUu8dkpIGCECEHb1/ZoQGPEjLcYSBSj7rg8QAVp4eYGJmkmT2p
PG1SxwJyQB+S2G2WnQsf3cQBiTVYGKYamFz69qlh8LzUb8kBHTxDDklTXD1/CngMH4OVr6w7blwf
Tjq+Pm6lmCotVd2J/WPSQh6RtDpHqep/kJ2iiSxU9f4cvamL/rfkuVDKL3/PMkzDsCi8XDxVfI/V
AsLsQnwWgdBRdHy//nvK7a0J02O80JCEWi6+cIiQlSEsqD+kkL2WHAtz07sIfI1ArQ/dTw+EsaRP
mRxaS8OEIGLCqoMfQFmXEc5y17xmFXKj+1mBA6zBpQqUf6pK6FiyGQ6giChUX2tdaCcWTKpfQuRr
2T3X19GDRYLMfmif7uXbbAEJKIyVMNWh8Cpo4PUd4iPkJa84JmluMWhPnj/jzqjdZ7fmQ8LgJqFo
TTWRpcV4pgROIf192/y5tCCmJ5tZdAhq2QEBl60an80PnNA+BQrz+VQqH324VNZuijvrCffnnqb/
gM5diMEiRtUk4JiXIgZHrvKNnu3FhgM3Bg6v0b5Gv3Tc2Ts6XRKoYkUKkYviNgG6bDjBeETA/Vc9
5vf7K8C2mPrY3enObmRtO9n3FSChso3C7l5IOYO0UbUfmcRST2+Kmq260UYfobfTzTXU1eoPt+Qo
aaNR57MVKE0AQ14GSsMR9hVYzX3LxlDbVCPU7xCp2wfvJ69LX4BEQ/dAvqQcpsGuEzEtFivmAa+f
xwOMOrK1B9lMwA6tJQEn7mCg1HfSTQST2qW6sfjMl6L4uniQ0s+8yT9kPqvk5qGhgtuA1CPVqqx9
n65dTpCe0s//QQx42NRnSxVJRz/lOnjGlps7ngea0yFslD/lvVZJfqwjYU8QQ1KFRhUPZC0durOv
EmYAAmPz+wBtNH6mJVkWxcm2ly+qQzYMWyoPgE05y6DIDhdVlL9wCSFbg65Hjea8vRyVTMvuTy2I
oyOSkVhZOsxA7xoUrIU7OezaE1jrcARjBGvi0B5/WYI6SdheBXqlHAJg3JcX6/jqdkeTvTeEdNpm
6iclyRXPaw9WdMjxMu0xXbyECwljAzy/hfc00oRS1CJXeEmhoNQcVxL1WY2USn4p5MqQR2pwXWaw
qgg4PSxTWVBPSUAFjJxmnNsTknSis2Xb7vvOUILKZVqxYG70sWDmpQHmTXZYpzsPn5lH3hiSGsJ8
wWJSJbOeJZOhFfBh0ICwKqhQItzwDm4Nz1O52n+j+eLP64qbUAzsA8LUSqGZtMgEuklzyr63nih8
MrJJ2chPxGX6/pEoN0pR9u8yccPcZ5IFMHKlbyHUZTKTzYY60au0RqVarM8Ag5WYGtDU64MG9mnx
ecer4YSwBYrIPgAssUgzRe8iwhCLP+ZhcihcKhkLpajPWeh31Y7t1YXqJK3T9CF2DpjRhBH9SKFz
fExW3+k4hmLa9vVYmH1bnAtqmuXuyuQ1YLbXSVipzN4hvRvFrD4dfoclCo21UdGpD9XDo9yOzefs
b62DXIgoCD3ISpp0YVYiSOCpBb/MjqoNx/VAznaEbppr2vKQ8rvP6Dah3AOX5bdX+qNp5C3ITKtG
QQAwwtZ9OECTeJ3m3gsTP5FIyB7+IC5lSAtJi1ZLDu5/tOvd3pRJbhwgvgNsQumeV06hm+P1TJcn
gVcV7AqSsSNvU4+GkPTn1XuZo4clowwlaXJRIClV+ThzL/kh96mHMxMIK8sZhlNnX64b0c/+864F
kMUzMQYPv/PFV8B29Z0vtsjMUgAt9oH0YlRPbkqgvvTrefwFyttpSscJvkoUOgiIZZI5BeZYzvsj
+UDU7SrYMq8ek7LJ9RoCCtmfdTYy4pwInvnZtY4jGg5MuG01f9ysuKqGpUbB1IImOjoEDWDBREtk
GDgp3MHRMpD59B4p78ZU/OQiwLqlXC0qAKoCHIUahUb9xXykvpFT2ctRwfVT3a0wgwBsMImvpq9Z
dtY9i8qYeH8PHhtvA5IbzL9ytYAuf97wwtPnH9M9BACn7ftC0jhedv2ADisT4Cw16FnEYaB0NtCz
4R84/kbqLDBCN9zQuTxGViiNNyIs6xwBytGljG5IoqzSi8d1XV1dGEb0a6bZ9/JUDQmgjgRY4ZwT
J1tA8RlDYgmS6l0M2MURt0z0nPd/uTuE9PqxDAy7rnDcqGI7uGIDrpB7FoAqAJG8+bCx/22qqChT
ZsoHaW6QgkFUOd9GolduYE0BgTHuYpQPnKhGz6a8CIi4ZkUKaCMTj2hYaC9Imgx2SWLNdvNbcb5V
TNR8JGUCW2Cl33aN7i09dM5Zd7nt2fxzd7RxHCPF6/9zVuFyJB9/pEGQrBZL/QW1AJg9JGhFQFuk
GWtMt+8wvkEGoEf3PjTJV3yD0DHbaKrJKHCcFYfD7ygHhWXJSkwSEi3x879vtinchu8fs7Wubn3d
PFA4SBmP5emoFFP3PR/LPPQQ7m5qwj7/9/8ZP+AnVIGEcGC5nSkjbhGgRQAeLNJjVzPB8YH9pXnA
c1Dv8bQUw+qV2r6NybHhxMXtOFATKU5bUt7RbjZsFgY+7Lj/HqPrcRXgWOdZvFbOfjxrvm4xCuxu
QNPZcQZz/7iLaqvDpZl70zGXgXbhO0so3P7PIemxQj+cl73nd/ygM9PboLAkIO7PtMhnNDtTiLL/
UZmSjIjGykoOSZpFaSi23jdsH3tT4eIwAceVrLOuWuw5DtovxKikie+TDcfYrVRERLqw13yaPFQm
WhChOZVev60qzbWJ3n0TWPTwdmaBQ67QMTX0koKPSYEHio/e9D5C1036zix3SP3W9AstiFirs7t9
1heq2dkKA1MCckBlK22pdDjDDIm/QpmMMxAyw24whSQppUXkNLZtAgANOGiMYf548UYt6DyoDXry
Ji9IkIvn9Yfk9dZGok+BbvBCXp9PN4OLUJm7i8T5YOdcr2/8L5rNZs2O1+uKAsi1oRB4X2njHuyE
wTPCiG5DkXu/IJ1k3SP7R4urLh4KC700pq+Abgh1HVkJBCCkUcKEQbZhNxyqbtc2taKxqvjHpihk
vwn2PuYxJlvGy3TJbZvpnNS9CnnuN85TCYv+mp9/KVgxus7VYsiWEXDYT6xyswd7Sk4eKpyWs7ft
DmZcM9qc5YsosRZNXdGL3o9KIR/rWx3Sg7DrOqNkgohiOv+vyaiyQgyJhHCY3dWmO+PNV9pszCC3
rboPrdb9KZ7SmuDdvQGCURAWs9QmgXq4aOgItFl4zpZZDDSZXejE5tIwZRtK6eRTya9l8ApLYtF0
Al7dCOWQODOmPY8fvg7fWjf4JjQrzTl3gIFD4z3cI3qkFqV5hV9LQ6wnbhKj1saIw98PPU+Hkz2P
6paNeXcKVmwXHIRCaLgQOAnz6WTaxKQoJOWIRbM3TbCCRrGzyiRzPjvMr4/7FM7vVl6hu3ouUeVo
aM2lpHxQkgJMMqluFg2+cNZwz2+hBS4EHW5koboLn9+VeGqCvDwZOnBBCJciL7NPwRFQpZZxqPPg
W3VH5DuZb7Rq1xEa0idTy2+kI5EK3W8tHesdUHkkS0vxWtU7gQB5rhK7YQ8Y0wxi9O3M3FiqjLlb
DnzfW9i3F6rpLgTebDoo3AKiON5jCHvs7OSbqUr5eZgeeHNJwDPG4YTKlJC/K+2Yy3DMDekgsvhS
Eg/8QHWG5oixehXC/H+nO39euQQU7c6Cuh/gGwVl3XWSJ/Fk7oKVXxiGVDf8ZhGwL+IP66uWrHOq
Ps74PVCOQdzYr+SOsyiRf9CS/kfb6stuWHjAgKHa7a9wdHj6hx1EplpjG523JwEr6i8Chba+0aDB
phPRuHrx6JCqNlZ0KghEbHVk9baMf5kGzJdB5wYZj1X4ubX5L+w+r+wqh0WLHjAIb5a8doZLHnHz
INL7NhKnQqWTWLRrtVYZi8kZBray9QpGXFJ77tRov0pfC1/4Kn/6lohGZlI+CKJ9jSOy4EtE5ato
OWvuDDNVBDTm7Ehkm4CW8JBQrvRhaRXeI0ZAeJjEBT4TzthWyIj6pC4EmGaUs49OfA0IOq1po13V
xr7dAy6z11H8YwvFsdqsgKslgAkBKx40iG1FZtIyceOnOJioM9AuShauuuZkKcasGMkPhu2J3yx2
2w+7pCtLxSNTJG1WNT86YUzgEeEFNULycCBC7M6BGl98smjSUlRJ6zReDhUQslI+JtHrovArHsfl
g9O/2r/10iUTyRYUBEHj/m7blWxxPIjGWMV4StXKLjLmuwtJGD7z07tsdHNxVBrS7y2DVOimf3kI
J4QJX/0+xp8HJNMREN4QoM0V+vJQNlB5Fb2oMSNVRcRTVKmTXlMOT97kOsZH2qMgzQ3pDCl3X9xC
cHy9Q3yzYj3tiqTHUawQDNddTxATIXkZKsXqO462sZvRs0pyhwwQhMQmvceIQKPC07JYcXHSdX90
fFwjGgFiDS8DQGZYxCXopbG5FRHtDk+UQumeJBLQZs7UGK67NL5Y5yo2JHFjL2EeybfBLhQgt5YH
4LT7KWCJlER5iOlb0qfyE+e4y+msv0rloT3nf0sJyWGAkjy1MZ4vr++euknG3X0Hc2hig/d4B/ou
+kYx1wA6iVxUPkDjJaOtyxjje8ynMfNMaRdBrDm9LPMhq8af2KbvMGpbovgzouC5DP0Mio9yPqzW
HWNaGkCEoBM6ICYeQ8NYhk4dLEqTOeyg1tXSTFtt6qOFc+DIfmdqkgHU19zb+O4M9NhkFjycjxOI
ZxMAf2Fftq0/BJoylzpuLFv2VBFHLd4WDd4Tma3mYaPfNlujf5gJu/omqMNiab4d6dAd5wkzU9xA
IdxTIKoPVnfRK33Au9mHmxXFToyjUyrVq+TNJ+aSTDjXBuKjz/1b1JBkU+VxLvLfj319YiHd4tsR
UAbeeDctgMaOa4MsuTuFHZ3ezO4t28LRzcaavB6D1QM36g0Dypw5BomXxkL/3icBt1lppFKnpPqx
41X/S99fqIT7IyIuVK5mCNCjWvmb6AmXIxztvu+8CUowgzN3lmVnNQD9Bms/A0mjEz+No+kObnfT
4QaxDU2Ih8UAfTnRGBsFMd3Dl3GfyXp56BVseXLojVGfXEjQ9P73WVgHbJrOeNK3XtOV5pyWCjjI
XykQuTtAn3hSAohGX6O64So/7Z58ds2e7PExtMwneVxn2ZECyhsEHwCnpCimhdZEfwebF+1kmgQr
RBAfheLFSzJojdCgSiXTcwKbbD4LnY/kvzyr1lm4snx2oW6gyg1mAZmZBLuqNz/ZK7qvjefQ0cfc
wLNqSebQe5MWDO65VAcEr6mjNQomYN3vtrlDFXT1p+1X0Bj/baMdxuGP1j0nGCcRIqEs3mi57z3G
wKwu8D0zj07nHudaMdr2Twskh66aTybqg5nkR14qhHiyybEOFFRmIhThOBPOtGU/TuFD7K2s+XfJ
qX4UcIBIf5xUoMxxPUJsr0gsOXaeNEmKgEHp9wa0pe7jspLhwemX/uklQiunJkGWy8C/q1KQVVqM
WvrFGgiZUNa89CgqyCvZzRnnG1rYeNzv/PnNVHZ5klLwSt9X9EcG+ht3yiWsgreVtSJORVedlTiB
g2hLJjo/n834oQ2KCwje3vFpI6UpnRTOGio1X81BpmpjQ7vxDzFVe17YXkGzFr/MG65DtMOrtdeO
cnpHYESc3B8xswufV8aoS7i+K/4RjLLLMV7e3b18eTKYZZ+hO/gTwaeAvHa+mmjyTTGG09/9frdg
mKJbw/4lGYmjIMti988kWHXIYzsFsu2/Z9uoInPhnQp/bxfvYtHHuP4zZ/RM7GNUnM31z0vaBERS
/UZ7b7u82BBdSsyMvK7H2yLVqutEaoyUAORfGeoipHhYN4eeoMOTX4c63jp0pELO69UG80QXJNd5
PY5zFY9z8SnIFrQLrtgyZEsYDadW2+wZlr2dyQ4Cvxdl5cPLc+0GkSLLPI9kP868vcZDdeLCTSRu
qYrdRszwWXDsUAUq4gT8N6Y25aGniL5Sim75hedLmAED73BkgTO8+ZIiEJK2ieyFQDTtSR/cacM1
V4vqpdQkk1/1wrng57hzhY0JoTOCpcC+xGS9NnozGkA97ZHQoDiDSUXXWlY66aPBnxag+Oi473IB
uGptQ8ZrYnX3oLwMWPWlzK+BxS+nPRAedqv1VUkc8/EVycKZqRAezFf7aRW/Wdf/kKsqljckniH7
AXcMuNaktlFoSsIAUepkOtKUIjta7DERM5U7JLfCVfEWnm3akjZRIeMHnMXxSH56T1Y7O9Vpvq7t
DzhiSceR2qHdD67MHUtgy0Wa2HXoA0cdG3j0KCudRqhBaxHOZwOEGr1WbtrLbwKH2h1K4OyYYCPa
j6nfPPDLdNt7o5fYwI4s+X9bbciNgjWOkO4Xi7GPwg7NfPKlHtsPuxHDzZ8R2J5h4K05+ayCLqTh
DjouOCTv9uBuTj45PwvJXjoizDFDfOgx8f/4B1Q09j91hxypPbqHL3Allx7Zj6cxxzs7dchmiVKc
me5ZHS+sRVLV7NlNxZ7BMJNw0RS/lSJngx4xFoPgwKrq4AnUAR565v6XW/4pb8FHpCZ2j24D5ma0
lVEn8SmaG49U/ChWXXHtlqAatMl+CVq0nZLyfTE5f88utEQCeiuErVC3m/N9KAF+edywo09i1b3p
9hYxCLivUKwHqfe0b7pA9JWzLiqcBsBqtyxAdoQ/eLGrszcbe3C1lH2c9gmUmgIjUDv3awnc+ern
OJyakgMDWixm+6QSZReSN0SqSsIC806hGa0Eo0FZRf0yK81aOABfb68MucErcySNQ1sxQ5OlDurT
tXUiGuluNyusf0rHu0HJGoEnfFQL8RkqVRGIrN9Rgxg0f0hKshsnxtKzNp7/WFPa2Ia0rC07WzvM
llgt0QawSqPS2V3IqDCYkPo5GUrO5GcU5fqdmE+GxsN04O7hw1IoOswfvDuIrlJ4MP2cIP8/KDmB
/RA3YHEZaU7bbCYiz3p30473KYYDQFfxqrGDW2u5NXe4jAAfYk3avrG4AIaodpYreWGMl7140Iav
ja34N6SFNCCKLUIBGv4wa5cSMVPPfdaLMq+XUS0kWlrHt7tHntwuEFp3aEkivTbAZGUXFbXTtBb4
+9Zsxn8MRJJ4gbJEpFCKIZLu5cEGbQxC2YqVjoPTdNQaeMYF421iTy/PcBYe2BDF/N5lAb8nf/bU
2t3XtcfAGR5/4uorOV2LShx0kCwUGrc03ZcWkDMizYmbCs8bfRRfCFHhh66JoH1Ie9uCO68sLNYr
QXkFTtfOovyfVfCFIqvS4V4sMJVPfyjrQ+jqPLVje/vODSqHfaityHmt5JjzLu4Cd7tzJVKBopat
F4bb9AZ/EuYWYp/L6lAukR+acKMuHuIWVa6QPMqcUhux1qHkfvvySJ+czsLQfGWd1oYMB/EMbfW3
D1M7R1njR41bJ2ZhDgsGYXvfP07D+iz8fUd5NRH60GWf0PnnfQSIhu8rz2HjWeoyKmEWbSaqtsn+
Cglr6n7ltKa5qUW4oVvq/zV46L1iku1uGCEwVYMyQSXLph2OEZyMi8w9HYgvKQ54g3huiNK9HXQM
tpHuqtJL6tXWgO8t1v2RWvXn4wkHwQB3PRWx8rU57qfMXGhR69L1anaR2A1/cQsBC9xHCZ3jBkqG
3jGDPL5FDZ7dJ5hO1jsgtshbKC+f69v/cl5UQQKSjD+JjrY3tk881Wnrgp2zymjvbNbwjzLWE2vd
E4tE/TA/U+iX5X1wBSxiaDYw9jdi/u44Poc0/bhpMeVyHJPYD9tjg1dWs/1deMMeLH219XVvmDvb
Oi4UGJUAJ9IFTjdeVE6zDs+n7Gz0kjvnNS5k91gr6HG8juOuyxouXhXMd2Bk4dwzt965D/sPI2B0
et0QSGpCx8tDTc1Fu0MDTiewl+6ie1VX5MjjYkdYgkeMmOI4xpyjnwrfMTuT+l6/DuMyKQ0uBiRs
j2B5kQkmDpu7+ypNCwyVENZFQTWvjYH07Imnf1bTrFBMzXF7/K8/UWsk0Me0JruoNtnZJxzmor7k
PQ5Z9MnCViZCBZuPHrUU2DKruM23sdW+VWio1SmIDKsnZLl9FlnYvFSXC8PE8sKbFuenzeJcRbFU
LaZcbhMgzykJydKRMUL4kC7rPHbpEiuUPRUY/IveETub5HxS/BtwN+h5fLxlEqeU9sXW8NefnqqE
+02l2rqTb3E23rBVKc7biULP4PnDmoJfzkU3/MfqJCzhEKA1sc+14NsemeINbwqUpB72sEvy3EDP
j6pVx7MbxnenlK7A5BwaBOz8IgOHyGiXqdWaSJDNLQiux7uazwyOX79ctYHDNZcVJHoSV0mStn+U
Ll51u/z1ouZerP/mpMfwc6v59yBz3oM/G4tJdxNCx0brmrT+k8yZIm+o0gL4NYUARPkl0k2YQgJE
rbJtjZtp4zo9duSIwCjeM7kHcN2AxxsOGUodIFwi3TesWkMlCtRdCeREAQwPSbKiXXn2d+7bnqQp
EXh//O5bOA+RxkTQVhbNr0bg/dZnClNd66Jah4i8sNvaymWamK7nOvLqZYfK6lfKrMRGhfWAvAzt
rz6nNpFsG6H5n9fWurXHFLys+8Zg21JZU/Qo5YWpvrxgYH9X+EHaWoXZ1542gzBtoCihguYe5B9b
KvK1Bl3b1XGANDAmYHKVOK6QphV8FRORXzHprYTFz8l+NDDdU58LO1AETAbXOJyCkHQhcsTKeZYH
YgXeAi3FZvrYLAzS6ndYR9iG4opVDaN8mxSEq1YVOpWQeCizcFpFLgEKPx5SDs9u9p0jj5pliWkQ
sbSfvi1tOQRdrDVnwOfVv8Y6VlFsRZkCYBq5xJo1hSwwXZKO1QsaQ91ugQ1LSqeo05xbPJbJNqF0
y2aZwAocd0ryOvG9eQGYA+tzpNgsrmKbCSiJjdt3pahoTU5bhwAXkubzyOJ5oNB+xKhjeAy2mWOs
ICHROBfHcVTAZb+0NNfuj2WafdWMXyc3u2XW7l6sguC72s0kybTrTAhig7c8YqhtWNC0M6V2orFL
f3Y/oipfmlvNABiidfBzI6+i8IriPw40vE2I8fDIxlip3aVrmXeTBFD2roDsHRYQ5meAw6R4XH09
cTC65eyvVDQB4tPhivqhfJfclgupku7Z8h8vGasLHJzrcxFTuTkyVWrs4tzrluYRFieEjRcKCB4r
VXiYGLNCke/ikt7jBYk008Y3ggsaBJTb+x/omQlqudrBs/mmcSBUOWoR1VdlQOmjXs/nO0RJse5y
4mEvju2YUMveO44gVNXNxQSLL2FL8dOIBTZYJAXAZookAeFcNkn0yM1sFOOiP756xUbaC66Ypnxx
Pruwtoj6kEE9Frz8BMD2zORuvZY8D7FDZ/yzUpBDXiLS9TDk2I+T6lCtc5veeWRbXPJwfpg6GVri
CVc3e44lgu8Qn54gGer/bHgpHiGawQqNS/n4GkLtYs8QZ7wuvtcrqNT2rGY67iUio3Nfz8ZT9+Ve
bqfSxIoESES+sjmXa8AAdWyMM7E7njRmgJsoh8KJQqnJN/nIvLqRSQEVcOK6FUzicEmygH7OQuz3
RE8r7yUKu2kK4alpYi+csUFL3zAjRvzV+s/z6ar69611FggRw3W+TBqIq5slSkCsX8RlOCG5Gy5r
/V83QqXtUv4qL4KUxPrJpr4JmwTxlSoaX6ioH+KlSYcAsCqFTsmG1ebVDv88+gZv32RBDpIngYlu
AN6wEWnD38DC7snZRxqIlLGTHLv9kXBAkO5vP3OfFY6x1GVgVpHVHch1qXEG25SQAN5pwTx+P+Va
8WlEsOZy5ttEXyzxe3Pu3uDp3R/8G9OT50ZinQPIiQ2OiUXCzWUIH8dLVwtnZ3hWqOh5YL3yx/3x
etXNyi92H5l/yCcAqKVI8DEskJh3j4aqoJ13Rv5K0lTllSbGGORNUjNKqHLHpJRi7y6T9C3h1uNV
NBL1D2OQ8GcUdumOTn2/qLVRCC14fRX/xKB5vtc+AgGnAI9tgJHqf5IIexReEYyHMeU0kQFg/9lR
Hw9Ihzd/Y1G/DkWkwIV+wiUFLLXFW+kdm/8pJfnEHFfzejrDJuBav7OiglrCYjv/M1YYVKWSvLAz
xyKFj90bvfERvftyAQiV/p6nVAQfqKbQDOiw/Qx2C6lbXwM0vBkHtj0hzNZ0UYHzzvC9YDI9eiKO
z5h1BPI8/iIJ8vEK4MKmEMVvM6cwAGrcZVLiFW85NFMdxnvYmOpNG2Cz0W3ldp2Pc73euk1brNaQ
fDzmP47MJ31MRecHCUB+UsJRwQpi+ovGr8orsqiziU474PHxFvAhV24zjMwzMYXr/vCXUpVGk3Ex
A2NFwRYYXpWZHE5Lpf4KJ7zsM8Ry+XmZhPv9bwgVSmBR0ILE7A18zofXH3NQq+1g7Pg4Xva3jJ+F
8kH46VJb9k9sXlyzaGJWLufVyl/nxoWjMUtVKNcWswQRvc4EJAuHvWXZgQm8/hKoMXbUNLv91h5L
6Cj3O8mK69UY9UMwfQUKplyjsNCMPUi34XF6yUhGKN0ZD3hHwYlmidEyPKn7O99Y8jJTXiaQ70AY
4vqqvvCu9GtNXPLiM1J6OEo9h1gW/QrYhM6w72qfk04SAGyfXkiJnYR8YbwBeU72Pq3vaHyy/YvI
AHZSHrchQ/TftDD6GWRqFDkR2MBYftM63Nu5Cpqtv40SR90eWtrCBuYzMpF4ckCg1nVFiKjNfOsO
IOEulM2iEOoUYOR5lCIveytFctmm+lqUfThmFjfzngKgNtydPST4kyiwUMgcLX2kY+kVMswYpcxU
t13thYTOPS6YaBnZM3EGAFEGVvotrfQUQzYEmozOW5MKTDHh+dXYHz64b7YQCRea8+i1WcrskDW+
EXgK4y5Sdj9v+I7Gx9cxrkQ/7dxArb7AOWoMv6AYHJCIWedS8k3kkSffQUH3u0xFDQXslzTgzatI
57lN40p284DhEKLuPrA7WXd02wKX1LiUBqEarbFi0hlXpD/DGjnvgHiQ5361i/thISFL+Jcdw2yF
2o8rjoGYi9kWEgkfOkkzWhiolIesPZXpuAmaeOr3qB4IvAE0a14uyZVXstmBd0Yy7nqLEZvTqRb7
dxhQnSXPJ1jzKCD7UwEmgTNn4etZ1nRkhkMDxV+fC0Y03y+kDFwh8sEZ0eU0RJUO30GSe1Tb8tPI
FDh6Z2Ll4gcgH8N2kaI9PDGpCbLLqt2YLJzxLvDjQWHh+Q0Et7aJ/GJaWenuSzXNIKWUe0/1OOs2
Ca9hLJug3iV2Y/kCgTzWsfbAWdu7zb4c2EeRQL9VS575IFktSlCWNP9C5aBJVRQnZ2fuNGWeSqxg
kbUXdEhEIcmmTS2zSIAXNDl/zVlEw0DcjCkBN00nMNKOwMySk7s42LTAtopLbAuj1XLrpFCEDHZp
ErGbofjkY+CGT6GO37mB+VCNtK5ukV4l/L40uZ+eD4QHiCPm1aWGNkRnWcLA1R4oqwyPoovVM/O1
85ohg5jwx5pPhaKNniMOLCWbOH628g1dVafEFPQPlVuIMNL49vC+gO7ZW3x3myxrup6x5x8e3/hO
k7eRWqN/YBXdYxKPm9ZtfszSAlv/exYYfmmgow9zucqFBaqEwkYDP3nJELGjpAmmAKBOm7ErYcCR
mESzwtB/RUSMr382I36SPmKXvqOjCztBEOEUlwuLNJt86ubfB0qPQbrRYt1SmRypUa+AVJRlicMk
//1htvvJYlJKCJ9wH1JSR39jBpxY0tEyw2vBLhrWnuuC5n67TLjsPy/ivOidcuoJMrQ+Wgp0tVss
XJRH6hkw6E+qz6qdWpAghAPKEreL1/27XXG9Opm+FXg6W+7WIXzWCUw3VguUULlaX/ys29oyNYmd
sSIychs5oH78PLwAKKOpYnGvn56YQq+Z9YQXq+r8mC1L5QhMya3w35aVX62w/eg0d2bEwUKlwBtO
xV3qnAQYeKAcFeLw14csEM9Ut9HQlQGMvU2AeDAn2jolH2aK1SROlY7FfVZivBBephChijrsKd+L
khXqqXhQnYr3yTMChmhKXwThYG2Q3ovaeS+PdwGYVU/Aw3wxZNLcLY2NWM8YjNS3dSaG3AKM0OAX
IZOWMHHn/CX/4DozCONENf9SFYQIsrJMraiwWgyOOkqYYskbzoLfK7jFGmjXbO95/csULMX9O+FI
OO3S3HU+vTWLGI76tn+PBrHSw2vgxPI/Lqw3WezQ7VophDSDVKmN+1hllRa4YveTv/UzZ4O671Ys
ogie2i3MAQxaZbh/mACzOgVVe5NeGCuuiG+LTfTdMncNcaPYgJ0LF3zVIbKg2uE0V6+JzyB8nZF1
bPzdfbWbpM85O9dBrzVOrNIg5y2Jfhtj2iXTi0In6qcEQ0/jO1W2nCW5jm2NHGpRfltpV9Mw/L34
JqsQ466UMreh8KuSgDr7/d9qxZw20zKtCO53KZfUCMvI83TkrF0+5tGOHv0WCh3vZQOkPtgycwpy
JKnu/yjEchM/rKLTHhs/t3Rm5tIQl1kF+GPePZAD6z7qzO3KMCrvuNkCDSTBBmCDFHJERAmB5I3q
hd9sFwbMVlUPPMw44EVMdWocMWcwKhz/1wDzpJEi+S1WxXyJjHxC+bIT+PwKMoIhdnsbqbD3WkzS
OIQ8CepBZ4PI97Ju1xWxEEvGZePYEj+bIfY4RVEIG8jUtFAjFyv42UMAtZD1NZ6pkr1F+pmLzBV3
4A2Tc43CiSCIwxY4KcWh9IAYKNg0DuwA3JEBQanEYsQ7ujI6lBwuo5rU0wJzRPQ4+c9S9PAWpG80
LeBTaEtZiU2G72TmsrVocsR+e/YAylspNPG5CvYZCMh+y7FLgoIsXKJfyXgFEtBYPwPr83F5zkzj
Ae0S3HOEBvAgh7K98QgQS0ZXPuCYm2ZRnDz+VxQcxL6SdWJTFL0DvIvDS+ewanvQIOnc69QU1FLo
XnQAD4OKuKxCL0oHJ1ETMaXUTPLKO5f5LoYY8az5o5XAvboNF+pUezq8Z++bdhRu2CIEUoLROlc6
YUloYZBRIen8e1oeyv1KbxUmh2DzaEe6RgSBL+DZH4+zJCOiDGn87fX7z88tSDpZcnQFDiCxARji
wSLC3Et6HDNZRvBrkQiG3IWbfYw0TyagBTPlYs5uJ0a9OhL/cVB4+HLUtN2U+IRe3CEZkPitwlcp
DDh6y0oQLWwgWsDHGrJmvqxKpaAxqSCk73mWtfM3slXw9XhfnCgrO2Q/Pfh65ckrcqIwnd5fiOIC
CHIlwZhGsd8OIc5r/Zt6rQnCicSHv1/YmQY7yN1BiobEwqDRk119TGZCWih49jt9pZZHMEUALPN1
Ewt/fSxnW9fst3aL+lV5DDMT9jGFBnfWZV+UiXdKXohs/JmTI56I+IGPr/XfU+4IikkrQCSQTHLJ
twQ6G3baay4Iz10ZQv7xvJyz7o0sy8vLWKht0oOM9lxKt6lhYNXe7iwoqr6H24M4dbw1yLk5TwHo
kZIwgAyen8GhmXy73G4DCd75g2cMcqEr97CVqGng25Fs7GQiTIYzRVsGAsmcYMzpgaAB5/eVWD4t
la5STWEjF84W62yI7w068j9IgXyh8cK6BZG1aMJsaMcZc0D5DUbvX+sDQukryjjefN+bsYa2bJD8
P/YlZYDSYUQzDzsMxNMzDdblfyvLuqYToiQkAl9x/oe0UnopQzlzyZ9+uPk9BFSaZ/mqnXNvvg50
WJdc2OQE/cH3NXVBOV+LhGeHbaDnyWSEqm2l0n4ElCj6+JN/rAnBBj9DBn3cFX35Z8SJ/tyWaeoQ
VHKzZhgFN0z4CU7DfcWRuBOuFOS5eXWiyNiIK3ZXAWIlPjva3xBJavqyX/jLDtXREByGli4UjYhw
2g5yvJuEeMN3cWBpHbXOxXqqWRg3+AjiSlnSXVYtG4Uf9x9BM8XviO30qn9jdWP1HeEKU8hDWus6
6c8lNCx6HW1yPfZeppAlct26nNnwTUNsXvEX3tiPE97JtcOjGY85nZ3fZECrqk2Ioa/aTSh/iOXf
aeaDWNSFztzLbXQi8RyWq6kBYA61m5m5n+XPonX1r3tv+HhvI0FiaYMh2sytYAiE0GGIXHmFcKQl
6Mknj5gPmA4797O1FmIjuTamFF52uQxAq1AuJhU0o+W1vvzoQw1SKrEhPVVqCJi+7Dh9ifZnX9Pg
hn4steW2jpAwyWx+VsVHG15qKhEaz7LoT0dUP/aO6E+88wti+f1MYSWIF67TJkkdFb9ePXMCAWYh
xTOlPxnh5/iCP0UQW+TptEnQFGov2dkpA7dWx6UdjTaJoatHK39G8cQNy/oIivPRfe5GtEDoeBuC
eCwvVw/9C5PfUj/fU+5rBQDpVmmcnUaHc2Q1QLNpY/7yNf0y+IiwRWMIIO13S8kWgQcXEKZDGsr5
hsYtGG3YWV8q4roKXuI8FqrroF8NLaveU2WWlt7TEJNxfk6bOuF894BlagJl6Z/F4CFvwPw+cKKS
DK1tOGe7e85TaYtBQ8aD40rgfMP3pxz0XQbwOLdBGDQN5jlyI/becno1kSV96gBkS5c9gJ/zBb8t
ISbCfvMavPcN6wK9CcuVvlpJLI+3WH4sgOZP2C2WU3NDVNqhDXyFafvjnwVs7k2knuVyoABl6Oan
ARCgN+3p0TV3HDWH7a1NBvff1R3NrZgZRfMFjuSRG4AiAUplZwxu+Xt/G3L9SLHHkMj7gx85YVYL
scSayB+7r7koQYssTWDRz/OpUvDuC7n1BE6Pi0n6vqmyqon2YijsEC3XyUWkWxj1xcKSCjEjpVbQ
kDSw4227vjY1qmLh3DwlceUv2vgtH/qn5+pkUBTCKhuKgKSCjRwJB/gLUCmJ2waZXYNB8Uh0xbhc
P1o2Qr5b4viCuYQpyvDWyyjA7DpleCGWEp5ojCpP2upsO4jATI+JxNW5TOPJH6DIBiJPEJuF4hlo
Xg5B/ftlXLqYKU3xLoAJmDHRnm/GqWFMdCqTclqGBY2dFcbwia9DB2MgIfOG9V3pEhI96sPD9Ok+
DpCGnoyjje+bKNG+QrE0ksd0RGgyvHLwtm74a5n5aUCAlD/ldy5j1ZvRJ9uVMI7JEg+kBmcfmrZK
Inx57ygofI2TiP/VTZC5lNeWVag3gQnlghSOkq1r7JRCYqWrlxN8qtXej5d8RBoOkUHWAWNarGCv
M3RmjVxq0QwJV6RhSi7H3/3oZTipRT3xBmEsQxSCTzVmqdzjznYOV7eV8cWEPDLWr43rW54eAFUH
nJjFmB4e90M/Mu9uCgHBvO1KXoe7T6nXPp/6YEa7YGfRlN3K5pBRcUVczm+8o/Jtg2VOfbagJPQY
t296b0rBi1z2ExJrRuE3r1/4gViQuh7BYEzOiRALr/t+WfHh6WrRDg4RIGQ71lnJVb33mdjsT1xR
yRU2K+E31Ols4ck5JI3OxxEZgTvkza3Yg+a/fp5P5B/wJzuFBeQcfNUbbNAKQQQs62BVtHLf649N
i4V+HG9t4fxDzf5K9DPHLRi2RFAQzpS6JvihbY4lVqQzcz11Z3dJntQkWsiltohF/7kc18eRjZQ9
pC/zKyemGNRJMR4QRb5uHMeTrnkjlbfY83pKiAb44Qw53J9mvXcNzDelHBUMErUKQEVl5wxFSnCj
+uLeWp8/CAm59dqQ5Wac2FV1ziRFAFIFOK4UMJIn+f1NlWZt3aYYtPgz7LLVAxoKe3PxPiIKKPU5
4Rwd6iDzLb3Yq9hqooFBzMfDUzpJO6JjeNtTiZMHnMm8OAxVf10OfgyHGi0gKIHpiSw80wmg2EHV
G2teDjg4KRjntFIBE0fR9D2CrP4Q+DSYE26J9QycU+8g15Kh1EW8uo3Dqzj1W3dBxx4gXboS0Pcf
2+9s7yhAbORnxL5Qak6Y39Su0qk2K7II3sgTVfPV+Y9n5Uu7DwDWjDc+72skuXXP0QROHM+4mroa
d9j6t59lOZ02OZeVeuq6lOmDmbaAxpzSOm+iypi6ndUVUc0YZNU3W65gIbt/Q3F2clcA42g0Yzy3
VALzIGcJY5tMhUXq9RzQCMPQipOqCURZR8+Vs8ISlf5AbLChu/BhpN/8PVopKA1OOm0U++tchGZC
9iqHgWma0//GEMV71ZlfVdK41pfCvLMQyskszg3o6V0J+dsDZIe0w1iaXuOD6/FUUApSQAnMtOT7
gAasyOQ564obCgF+DNTuhCa1eTfmqfZ5t1pMcrRtiE3HLgqKVui+utoGTTRzeaRaepoHECVXK3Nl
Ksl6uZdkYAWVDGWMctOcPkW0UR4Sw0M5v6ymHL91NTDCSo3NkgbftZO0vaniQpJHf6hfjAoSTaZg
BFvHI2S0vjUgLnK/ARPIufeZbR2feV7h47l5u8uEXS2LYxASTv/LQqpXH4/doFrbcwKV9j3QhiF2
LfqSINEbOc8ZQw0Tk6ur9tzSHpoOxXR1Gqd4N7GD7ObIfryn5cnp/ST37TjNIZQanKWk1sFpLLd3
nPxLHHTxkAEPDFg2W90oT3RzsMV5w+pTcGouWIxHsIARXiO9N4Z7uMDT8a631TCEjBVcQ03apJub
R7rM8Sfs+24sRX9inxU1E/yJkHfTBuARHxKPouDxQlQM5kXy3d6GIcAICqM0YXoLX+tiUHdiP61b
9TfL0Q3e9YHyV2b5YAozLSciY0YThDaHA9QUWMlMBWUEtz2I+wldWmxvSP33Sv+N43LxTpmxpV4i
1LqzhWOsHZ+mh7/zmP3blKwYxEOyU2aTPuRixNlLab7Kaxomry3GWmgsl8Nz2lqMnH+WMT5F4Im8
VfZW6G+x5PPCEJ80OTHW4fIMWULjLpZSEDez8kPSUxs7orX1+FTtCnyilKPqYRWLzzyAz8CnDNUX
kx8GljhpVXoTtHQ3lusSjKsAI4zrozODd3+xEvdC28Ue4nGL0OXZ1P9SriPCgpcWn7eSh6uO2Z8G
ga3SO4XP87jw4wMag2YvzvGE9bmw5wBHXUighsGCay6jGUC+HyUWmGiJKZ/znpN2/1iFXaVcAX6A
JvYXd6ualpKOE24B8YFgXBLl8b/AergiVHzR50Xt+UwFH0fBWYXIgxgU6BcieDGAHxwLEclCMjPE
g8O4hoPREwwCkEz9lQJDRGNNjsSvbpgIshGbZX1E2j1wA5PboYyYBxwmbtgXHb+Mpy5b5L7Wzh3h
wizO+iUQLpv7IvH9EPoeKUFgbP3nuVEbhVDApyF8lf3bkUgFMO7uXnUpwZWhC/k+HCCCbWPdeHBR
Gw3qXszKEKA+GN/6NXIHBlTC1gSBX1TNcLs+Svw8a0nIyXjQQAhF30/Mkke5shSJguEXZErMaxZI
6BYkYP+HmIB+Qu8LAp5WIWS4m2UDB0rK4Lly4aZ26041z7U6XFawp1YXfjyhS5MteX7G0gBFy78Y
azNHKAdpjSMEzEJgJN+OSuB336jqYLaooe8h9FTjR8ssYsjo3DNceAmULE9bbsjhdNGy8cCFO3eB
dR4PJ7KqA0C9uJiIO3RydYx33n02xMF2WvwbK/9I/KNE4W2J0ooXKLE5+h8WHW4oFFEQbCGuhcjT
ZMSf0GeezEamsQsAj1assQRoWcsvzgAX/qArqXNdTgCzDtUVCAoCxo4r8fQucTbPjjweqlqa5hcZ
WJ4qIoOuFxYC/aL59sSkhk63RLtkwEbuiiUCRVVadzONIB3c6cvP6MqDEtPi8LNR46eACEwtMsge
FxhcD8LWeDFJsE6eWAXZslDLBWG2k8VlClOx0S4N2FZRvzqYnNixnfIztZbuIPCameiozClI2oLT
SxyK9GhQ5740L7ahE5QjwaVnSpqyV+QnUCXTlGSQT60a/2jVVLts15VQW0L9qrB20nzPxvhLXJsj
biBoPZ1twHaPIHqM/gAhrP72kxxAfIgkxuHoKM6k8Zab5zum6bt6kWKmx/o07zeWvwQNws8ZBazZ
r9wEOiV9MW7QsS6cNIoKaVDwO8sn6i3HlYpxF3CRTXiMXDzV1m58MLLG4KOTPbHVSO1p7mBvAupa
lAbYz0EhaLtm7U6PuTL9VTYsRnRtkEReVED7vK1VK3yp7Zg9+By/Kvzzm0rQqF1HJP9HNF6Adqf3
WqcjPhHN6ibz5rK0ln4q8Ibq5eHkSKKYhBSlqAmY6emxvXo72wA2yjOplhSuWOG5smYn9TFFnwPy
IED0sutTyX5SEAm+S9uyWbKydIWdQwWuJQnbgL3PnnLi5CL9EY5gs74kj2yuIsbmXkjgkoiDNriZ
gm4zrCG+hcjm1ITLpAixmRA1Q22MHKKZtY+gcf9C5FGov9WR8E1kSpPCfFYUxbR4MXXwAW0vX1vx
acaTB4rZkWZktmxDedcwo9NULmPXs2vj3F+AtsATs0ZCRDWmQmj6T+QxzKFNvAqQD1stL6v1Zgwz
PinaQiKvoGN/90t/IAslSG+z7INxkq/Dn0SYaZY4MdfZzO0MmXD9mVnVPjKCVQ5gYnhdi58pAI90
ekC8A+hw6okZyT+11yFez8sR7cAm63INZQ9S7gQ7pNelQR97PXcBNhdR5/6kDbe96Xpc6ySVk8o/
Wo7OtnJeiqQ8l6m3YCHNFggOLJ5goXqNU01T77DX4rqUj/a6YzWV/NmhU6Lm0j/fZN9mR1SqDw/L
wMoAB0VWCuwfKG70L6K/QAFOuBRIsB3CA1kRc//4XOgP2O4ChY3FxlQmY01itpr8OY50u3U3pzTl
lrM/0yXFERJix3qsDwk1+OiLuz/o/QOAG3YpJEQaM+AeyzPNydlcGQ9m50J6aGFe+bQNGHxST+G4
+3Enncbo+nM1jF5rMwsp4r1/7PLgwdpEB4WzS8Wws+zuKEEHXwEU7YpExBj0/GbXIq8o83x7/sK1
I+3M8Th3y0osmGwKQ6c0Un4PYzUTESpnznugUnupa+HZIKnUwBjo7Zbej+BaU1DjZfG14T1jmEvK
D7ZoeFuFyWADzf9t71N6afq9sK2lWSZqGNj2wNKfcynWRyMfmuvF6cZ0S4uIYhI2P03qVePnWTYP
aeWSQLYbd4mELEqnBVLtn1Rs1ZUUotdGJA9ZYBQbcragtfYJyebV/UtV/BQwOwi/58VStH0lky6x
4M+SymFdFtP2MVS4O91+cu7YEwZLTqZ1gHGCji05sa7joVMjjhJH6NOJMXcY1ZamU3kGmOwCGKNs
CJJlgH1oNo9bdUPzPUl6KtRJ/foO6QrgUx0C/HMrdp54ASpEOwMGnc81puZS1RpfQqDR1VktNesR
QbJrGO8+cUFG4vREGaEx+wxS6U7BDFOG9gRsQ4qFCiOPgQmem/TW4SdgDesi7BICH04VXSB7Jvqz
RgU2+elwZxkWtaaIFxEsrceoiNBodC8hK2TY4OmVqR404LNxBgClptSf4nXRmbu1bTQjS8rpM8dJ
vot/F7u6njDt+8e9Y3DmULTRUP9rLXdYlIGaVzrDo/miU50uMNUxWdCjlkLNgrZ+e8kuFNBWYvo5
j8hCq/kLNZsW/rTRLTyRQwt7GQTnLotpsHC97jbftSaz5jq1GwMXw1b6qWrf5hWt9/g9SAFpXxZJ
tWUAwR9Qn2mh3A4BBcuwazi3NeVFb2fNf3ZF+aLXFPuQuax7lkG8VoIRJ7Gnw13gno/HBzmXfhbF
6iQio6DLoNGmSzx+FRSwTtR9ACz0YVmSl7xBudykPxaEoOMR5qp8OWuUIoNkygQjdSemITjnFZ2L
PdMLMoQ6i5RM3fzBSHshD/gnYoNj5CkYnjW94nwUOIGw5MZLqQv1OgbCvnorkoN69RcY/SuAjXGW
bEClcanzwxFkgsJwCCrRKTkDjL/GdY/t4V9z6dN+9ymuyPHrckwR1gmA2A+oI8C1HaQntj2PUylq
ebDEjrrXfR3bMMk7dfMkZN6Qi1fWdRvFQM3euCpTwFvFRfUZv6R5nYx9pZqKAeSBDn9i6asBb5gX
R3ttkfBGJvKqIvrosSJuwsmCNU+M3ljFymj/shRHgOqZ/ogfhTDOHCkcC8GHMnyEWDHjPDeiSQ9H
wTsTZqfI2weEEhV7ufXntqzjQP5WeREx/5xGMzTxhDXBkQ5TLH0utB0iAjznyReKxI3kggEb92Af
T72JDbrEDBsF6vinlVpwrse1SQRr8QVKeuTe1SNSw9R9vZVslENZSpGKcinyMZHjslUiGcW4pDMQ
ZoclQHhktGjifnOLyOB0kCZ6DJZbpFWUSg7OlJyf3DizsptkWLqxSlY9GZJy0vYQvogAGh6MzrH/
2+2juPZ+t63ep6ZDBDPWXmBaSXWn29RbD0O+kP24U0f3d0UzofqlHOxjow8f83BqJjguBxp9TBmD
IwxFn8VlZNTi9yZT44PrpmJZfjq7PD6f2xK6chWq0TzJ7OBX1BefPcOB/b2Bos7TtdR9vUepr335
ol9takHzIjeRlwiggExolQ/IQ+0B5EhUp90KyJ9HaMvGWCuo5r878spT99vwr3RIynKPwsOUZpxZ
1Eca7zunlrFr3TkMbEGytkWFK8RS1HFHVMD2JsuQqEifsxiYvMofTTVqYYqlBib4rikjVYB/BjhD
s0PkOc4pRezvgQ6kwP4bHdn4OGvw21nt4wW73jOmv/fPdYIinigMLw2Kib6Q61l6teNtG/E6GhEy
0asU+uQtLjeIkrp2cBMjRSo5gq9HZAyPLMz6QuBNC9k0PqTZC8wosktsjFJe7qfOGmsYQ9nmzIF2
uq6uronwuG456h2rZ44uy7THYr5VGmOAH69VbafBYzaJVfnbi2d65CNypX/zQ2nYbkD6ZyS05xt+
ZUDQ4hbB1EY6gHuDEFvko5k+2/rnlx3i6+udCZEw8REfOoXHIqP2vqP5Zr8ouGcFZcgqhosTxMzg
08RFYz7hiGSGbcxbCuk7ucxQEqq5ypVDkMscF3B9Ek0DtZPuQ9J//kYG/eGsDp5bN7IPGh71VjIi
JXAa8+6Cj9CnZjcJWxFCUv8lqq7+fwOFkFnC+gc1cJob+YBv/345RdSoYq7MXO9HjaszD8ZSSxnD
8Ug4GXEo6JGQ187Pz26J5b/t5NPYNR4smdCVT1TYIQErp1NdtlV6ngMH9q6RB0g5crJuHBFvEwdW
7rqrn1eqzQUzfbhAZDbAPVY0AcW3dnyMIJ3e6wWehAFg85YguzL+aZMk5vXNX+U+ADB6yiKE0lIa
BDpVBHCsEfjILOusHldcT36ZOCybFuL6/4pDzP3SrSaQko6rVLojYNFZcwdC7YSA/zFKjSXW5M9R
5G03qfPe0o/1mTHZvsnS9q1fq6k=
`protect end_protected
