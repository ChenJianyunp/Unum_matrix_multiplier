`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q9SNy/V8jztMyq4C1WWJ0vyeADMSOyppnBiKwMmuS8wV7UCwEQQw1F1grJXhMiL7nLeDSj1BxB+a
yiTdDBQBFAunzZkisZc3aSIC6fjUaFPA1ez4lgZdzp/3GFwQfOxIJr9DfEqLyp34lpxT6YbOuwGx
DrzJWFZXZMWNRSzbw+WKPRgX8XCw236/IFb40nvAxpYGHLqiImN1vuR35hCmLfgvGX9Ycx5mSWVu
7IqzHHdD5lZ8xEfbVGAX4jcesKilwx2Q2vGx4vpfbYuziZHFENBqhtNJXxlYO/vBhnsQqhsfxqHQ
wA4GocBjl2iGWeLQuPlu+VSziOD0ylYu8nabbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 138768)
`protect data_block
tk0haca7+iuXB0sWUwTJW40aBPMvgb6+8U+Oiowh3jeMPkc53oAmi5+MfoMy9tQMPhG/qp8c5pXm
yb0QA7d2sjitFUXi3YRt8lsvg9XB1VaPpYlE7nvyN7cvxQXIJM3bHFyzhG4Sd9OQa+LH7H1aHTOh
qHU592qtaNa7GLGarnqnEm8QhPoEvkZNUfqnLmNEJjQXougI6eMoBHBD6OuDy5kr9ZznB3onw5k9
QFvLkolN3egnM0BIKbCrj0V9HuXmluOFzpPbVnVSRQP/LiDDFr7nrrUcknE1KOJyQyILOIZi16JK
TttwkowDCbXpnJ/d3aK7fy5oPmuO0Q9aR2Jrqdc6GCugulQmw/R5FJevwYAm6AJ/qrKYwIMiuPBO
8ouCDswGoZLlyrL2ySO7eb/vQsXeQtsMdDYaRtNBGKuGlyIaguQ/LHE0XV8irRDOwr5yTT+FvNAW
nrUZ7lfrrHCAreS5ti0v7SGmvVdLkRzCXxElvLvtqfzRl1ADo+Fu/i2/W9jbz53uAadeEXfCYaFF
+jhlRr1c7bo2xhKcUCGqI1bcUn9B0hjDQ1BajyIxB9WPTIXFXlFm4RSc8ChOApg3ogXpBupHzM2f
b8ky4nIWIM1tCzrOEosCW6qBrECAavGTI27QJCLjkZSeFs4PRypphIirRwe6HlZo277khIAkR/CU
R3bQZc0/v9jv0Zr85/rmV1Tobnl7aZodNkM+395gJ1O+FhtUABY46SWC3hpQqws5vN65fmupZd/N
T01+63uw/8wfqiy4aXBRZXuez6wDOdihBbaLi5zb2fLP/HMZlG5GBMHzR2i2np6vN9x9Bo8aDGgf
Md8xs7pzKtXpoR6HjowfzJ5UnBNHEOBaY+0lEd+E75kSgPb9Z2ZujQRnVjGyncjkD7GBOYFSBVs4
R7F5wTSLJWIY98GG5bbAPa6qPsT5ZVjpV+48xh8PfKkmjkj8sanfWEV3ajgs+ZA9vA8L+NR4khBM
jrEXCxjVpm/H91xxzNlK0l6eAyMSapJ7N7SdyhzmkO3Os66tUBg/2UwzAS0uFab2wZOFMi+bMWbA
CJPNO/mHMJkvnRxm0SNrMnHw/dYOwL7pt1QlAw5USHEEawgvzquH5HqUw8CpDKI2tZu5fwS/9pGK
4cS2qouxiWk0rKZ6UDXe3/PcXUHoJMe6ccltkSTXRKkXuf7JmzCoUwvh31gtGAbd6s8TGHijy+v3
3DfzJg8CEmhUO8l/OcrDRLylx3tffmnBjRk7sR4DmcBRhWmrBcl+jEF+LPhzlUc/j0K+CDI4xhiN
5+uywXywyQLPIJkogX6GEYBkUnnBDH6xmmojotZRAn3+2ioZH/nMjRthV+5q0Nm2TLM07At2QE+g
0TCAE++uX0Ukd9HgMYtVPK/cTIrLjeAsqHcJA8uubf2/1vwJLmCC04AT3p7viojbQQRHmR8oJcIm
DrTWgRlPqJE0w6dW82r8mCzwsy2mN92Kpn2vFWcY6puDZcqTIg4iznp4X01qXsmA1FIDDcGfSly2
FGBMiQJpdehG+Zw/kPyRqhhsMXYOS6oqT6GZyJCdAZLwBiYYRmXthKADTwQ2XINrQl4VwKfuhrjt
xAOiYa8yocBd+fQx1EKFBkFPHSYa8Fad8bbOzD7pJxEjuH+Uqz2YBX7DVDXvAP9JDiQJGkodoO/9
U+WyB+LDDI/s9VPFAibFLJ8dJRIFqZOpvpQVRwqfDHD8Xu5VwS245T1V9k1Z3ziTXKEY8Zs8Z3zy
MLGfn3GHFqvVE+JASDt57oKlj+zxkYOnpuxFPLXCVf1EcJmXXzpACW0ccv1zErRyDTCyEb/tzIe6
pHCzP/oGrH1D4Dq0M6gASkCVod28WtEWhYGKX5Hd4qJThO4VsldY/8fAbSRsNu0uvDj1IfRWggXN
iHnjvxNbXCUHPW/qn3khc1R5Qq3Zd/si7PNuBTWXYdA//bezJVjHNON+rTXb9hcTHSAoS1PUGZiH
gNYYugaBPuz/ZHgVvIdZm4BYTtMOcrO/W6gUz6eYiQ8/Zf4tP+QrOMzXiZ0Ij4klbRc1VslvCCqe
n1j5sdIsX+oCH2mBlxAjMBKxHQPc1hP6jpJk0S4Iy9c886w34MPVqWO3I8y41SXpPFWPX2ADX76v
MDykoBXsVQHZYkzhe6xT0FZ1SoIrU62pBqR8n4fBbui01j/tnjwYwmm55/bdjTkM0CJtYG6G8HhK
MCC4VZZUw54GlJVZnsU4ZK2HhZe+zdDy7piGb7qU63WsDnw3NiuXASrmJCW4lGQekiYzOZfZsPLl
KY9HdAuHPM728kc5ZrqN2g2Zdyzwd17p04ndMV/RzHnQgb0rUjiDiS57VqtmE1Y1j99cOQkoUFS5
aJM95qheLRlD2A6qAl1lOmpMVlSkfMoDAu7ZZGNk9qF7LfBcYAo2nf6PX+3sUl6EKCWymcdmH2SW
u2eVN3FIdQcOzSg+/4O3pehP6GGGj8U18QIEIXE/mQbo0Blw4pFO2DTFfTy9Ai+0JcbPIinKPOoh
dmMFMKD23GbMj0c0zLY4pihUMGrhbfII2+zjN+112fjSn75ecqIr5q88e4Q+5gfcnoNh4SIExquK
u6Uuf1IiDLUgd8SYnyCuqZqOT4+7OsDEXXNhR0jDuvCHi11EGeJnNs0KLrlVw5bgvmTWUJJX5Lux
knHMox6PUVsD8uw5Rrwhb3kUPnwfOSkLLY/lKqHGRo3MckB9a6AnSbaf5+5r03LvSG5GwSnoeNHb
oERJatZl8A4mDPiLLrJd/ZlaEort29yFUi/Ol3uF38dnb0YmhK+jH7hBIW/hW6Rrm74j1ZD5XhQ/
u7uPRdzOp4TPsC8Xn3vzW9yIRyVjVWqRxp9n2iyl9hgxEt5X/6vLer6qp7P5hbeBXkQwGfLPOWzk
a7cs+fdP5DF1JyWd7LBWY96zJkqhuZxg+O6z4j+dzBz3iikVUw/IiroetuSeSqW7+VBmzrsWpjfi
CD3FD7/HnrftlVjDhZFUl62xvckHpDzbjUT4GilzmzPIh+MQC063u3ts2o9lLdycekMIKvu9vsO2
NzW35YRrjPCcY6NX0p9UMeVltDpFEJM+yhz6QLqMcyvDhbU0ISadNC1YekFzSnZJa3geUgPtSxqL
uerBn3F3AZ1hCYZoyO0DMFO7X6D3lRoOheVHMfh1t01kk7kEUxAq+rwseru5ocEXdXB4wwGs02Tp
9x6D9cnTk/s0R3u6i9x2hP9h9xVUOEvfygXhredo597QHC4xtHtb8k7uk1v71FcvLZ+ThZsg8B/i
JHkiXJTnJ0u5Kp63XfS/r9frzrVPYpHQ8gZXE/GwcGFqoJhpsQw2eTucdkL3oek+3KwD/bdrQ8NJ
zjh4mVMbb3nyKMYYP3cwm1b4eHAhKr7TBhON9ttVn4GDbE04ppkFuxkfjKYCwvoCDmNQ28ijDsB8
+xBatPlXhAllZCShisiN+qTowboehdBHODAkN8LrLKMqeJ3B790AFcMhF1fGqeIcUReiQUKnNtdg
eV6lz5alqY5HNbckZiW6zCoiwpPaIpH7MDZy3jN7NcSCZzARsuzyEfiS93ToF3gcouItQTNDDycp
TNb43AU5J2hbcuSLFT0SyXOGtKhhTXIM1J94NMjhgIuomnMScySTsOmsk2DNxhOEGNVIab4M6rx/
7QkId1JoBlCipCVvLSldEsSLQQsKTgQbeALjFzSOHFGleilYC6Vdo8hkiRqt0vOl0kjyF/mqqvK3
KL7S9f/O0mODJ3IPh6RK7paBnuSkOGb/YuVigJHnKSBFFIut+ZcHR2OyahZ2FAZUXw6AenOt36rw
mcJO8BarPQZv6bwSx/T7AIWj6U8Ggf+vQWZzWz7yR03+b6UDOOpfjRjfWAxeGaWfl1Wr2/LwyUv5
l/mz+xzBzg3BvOAQpfdTwqTMnl3WXD2l6RyQmRWVS3uJEl9x6WngyGaMH5+Iv+ZL6DNM17xm3a0/
K20xTniGMGdV+m7h4KeVRjxK6+EHSYo7bGislyqRkOCVaX4gTCtQGqpV+U9Re3Ioc82WS90417bU
IbGrvyh1r33ornrRMFyiFy63AE29AELyhuPrJLvQpAgiSYam73+IHmYKEnRtNassTxVPPxvcIK3j
pje/HPzWBN9lSQN3D2+E0+6OUWJz8/5KEWrl03OM8rrZq2HMO37H2FJ5w5g6OKmeRQRzmtkl3I6D
l14DCUj840yzPXzoehO0jKnlnHoynj4DvcgyMs19qclo8UEK+N+u2rqy8lfBRlrnOfIVuOoMTae7
cWGxsNlYhy62DTCe4rbLt9MFi6nTySllrJddyfwttawfauDHKFO1CSB5f0ckW3VGM5c8AXbORyRY
oQewBhTs39YPvM+QObQCEb4U14b2y5yPZEGBnd5EtPqxLIQhV3lo24gM5WV6w9knPZLbhzuPnjtS
0g9lLHafjEz5ASKVqW1kLoXhgHl0xQB6i7IpsFIy/XoWdmXL6Mqk6TgSvd5RxH8OAvtC9F8Gh8Dp
1q9JnkXF1jU0Q20NT/yZ8JYE24dPayD5x17yNJsNZ+qW6BHo71ULTNntXJU2UjC3cytjmYseXWLk
uF3YekcdHyk0/AjoWhJlec7HU66rx32BoFuonsFdfoD+mYg82mheNI5RmyRQCn8KWADnfj0diWeB
ihRptbfGcsvA1sdud2auUhDtMj+7tONZlbz5V/CEd9UPZC0ce7U3FDssQ5uElNx2kaGUhLPSkgzN
VRgtDtGx18/4+t6Iyg0O8LAwdLZS2n3B1DeRbpqekrcVKAtf71u8ygt7xGl50UBMmnYHzRy1bING
xGOJfSI3cH3CZq9C1F9kzLLn9XvX6GT1s0j8JXzqVJbJhLOc6iFhpGrKja+5A8eG5OcsbWPLR+6C
XF6Kj2oIYgEi6C3wmgWEsWLi7Y5/07kKyKfxJ+VPKwG+UiGztxzrafRMvK3RfQHFABC6wh/Ewm47
ek6KVT9TlRma6VYatQEwVoidClBoqWlzz0j7N4ZCMscXjkpOa2nBUoMDgF7Lt1b3/9OAWaJBPrI/
jHKn/oh67rZe4RIb61AfXjicA7pfJkfNOM3ILCIGprwv3Uytyx3F2UKhCGNCV8E1keqeJCyox+oB
j7qWMerpT10mfiSMoevakQocixA36HPbbARWg6vWRRrv5bzX0SSg15Q0WunqbGPAvSmexxysQrJw
q0WsbUic2fWLnvQ8m37RMnCqu3OG7u6n6DQX29eFGD7eEgEO7fDrJ4KBq7ZZ84+8kGvUt8Vs+84n
oeB3cHAlYq8sxDEsKkTsZGDuvt5e0aIDD9BftXHcOQ6/2OlN4c/ZkTWdRjXGV/emFIh0YKVRr9lM
+lsTEnnmSia5nxjeESlwOmfm4S9kJFhmeVeERaJaVFKDpNk//HSEnencmBnmxNvtZZbM7vpJg5a3
ty8V0/Jia0aZ64/VLtona70pWfhNeJIDArfy6tz88qbaVwNdxB3jcwfJHvSjtDse1e0a197MS7Xo
JrTjhp2ASMymNHObaMu52tW36LeOeahPTGGeu7DpbQmr5XwtBsiicyVa6u/Dyp4Lkk/3qRFGelgn
oSYI/N4vU0uQBCW1cmGzOVJbDQJxzQ13xHijY7fPodwqiDD2yJdYCWur6VMay2x3vGPLjKmiAY0w
FxEglEFwKX2f3p0MxPPs/vWIbFH0HJyngWeH4AVS6nHxN13mo1WbjUZ0H5C5pMU7nq03DPBgYMpf
BMgGTOsOVEUbILvOyHbUf8siDgNgZ3qw0NFuHaXNz4+RphhUwhoOFUUlavpLU99pEWzcTXEB4+iM
10mYQjQJUMP5sB/UUEHtj3q08GwTlhY/yEVmMVcKEiZRR59sczyGqTQVlaLxQbcYzwyMkBSnYAE+
QmfOOb+Harn22bWXnvdA8C0hHMDqV1Th97p/rmUK/K6ndh9WqWHprc/aJArN5rBpNv+wpv91/5Bc
eShIfEcax/Oez8bE9USkTDzAIMnig2Rsk7hUK3v0prDx8TEXNR/+fGQ2Qtsy1GmX2t4L5FuhqQLb
nKpHKasKlBe5953lMBYiWGWCLa1kP9xhcKg+l9UB2MowjCAbIhJvQVuQmHzFiqewzwLFNYjeFECS
ha/VVhyAroWYboNtHiQ8yqSU4soYCqpECoxpvGsm/KC57B98xv+TDPXtpB3yjPsdKClIv6bhy8WA
GUIysT4M1y28+zDa7YlBZBQawtcDFrTWnO8V8jZKUrVbARFgXtG0iImB52TsHFg1o7bEbDMBpg0S
BRMHMU4PpvHcOJ980aRhb7J9dZjNg6Jmu/JRZ4ZXdGiZriV7jxLIw2Yp8YDBy6Cg8oRkPVtX0IvF
hjjyWGZ2X58vvdrcn5sUAVfvB2rtLb95CGsSEUh/1mD++44lTGdQ+YPRcD+ZU4S1mUHH6a/+utKs
iyzFslT313ZuxFXuR5euIyIG10yy7WoQ7DdWjJrKYtbnpXU4YiBBqceGbCKLQBWovhEbOVoc9iOn
J4nyNFw1FiQVwBL2sgWCR1qkSqL7WzAhVyM5KAIeLX3ufJ4MR3+yL5WIujuv6m+b7VYvFwHlDclD
E2w3Cq1HDFv4R4z15WmShHEtjaXVX2NMRPTt48vXjC2HdUdGimO8keLQFjstD2CWtfaRYDCst+pP
iQKsZkpAS6RZSCbUAC6p+K3IDj0vBynCkVMaKCgxr4KCu2t3pVnfxLPVn0Ow43jAysmDpt/9WP3D
ikCPWG9PVB4/ErdjG9ldnQCmOTqaMninNZ/I+6Ykj2xn6I9FuQPzKjMS1ajk98Lyo4yhsrz5n4n9
ybn6IR/2mbcOogVBz3FDQvhsry8OPXD0Un3iMZ4ZK1aWiaxuJmx5k1sfWbmG5smd7E/4r52L9dmp
ZSBjQ+MnoD0W8/dZjxh3cUfp13+mavjtka5CbkamBUskqRVtBmUicRG6ZH0B+WqEa6JwO3JGB6bj
X3GrI+sLvxKKObxiNCoOFu5Y6vvd4fWy68i3PR+eWkn8N/95kflFqAPYaNNIQxWRIU3i3Vr9Avrv
/mnAyekhJBinNi300H95vTXYYZVW6dWE+bwp6xFfQNLU3bGRSyxdsunBgAeoKbX16dVCJBJlpbVe
FxnRaXV5weSRnSdAKNkL4nJ6I6QE4iXuCMVLK4luhQdPJCFdt4jLfeHux1Yfxu5DI+I2YhltJ1/K
RRwhMrYYaHkmtmkUaEEWd2TlznEoJmKQrYSEFxdFFhpkH3MU7POvyZ2xVzrDFf7fHPcAec5W2ntT
1j82MkuSDQEzb02g500we1nk3q5L+BHkQzQ+gtrNErlBepr+rupg2zPXxQy2cxHt5ZeFn+ClVUC5
eVMZokx1va4wE/yX4VbyZdNrnE0WFgaSKfSDxq2MENU3Q9NQ/jgdPav9wDD9f/HmpNLzO5qU2OHg
8+uYyxf3r0J+4KxQjo6LYhOkYYe7qG6rMp7UzAO6MfGSi11scAeOKw+851KSMayc+PBhm8perds/
DqxXcF2bH0sOK/+ICxjRT/kGUw4+711w2nY23YJWc8YVUKEuLZp7L8wcfWK2WnaOgBL2ajbeM5m2
+g3IjPZD7vLmxxrAAsiM3JWS2BuN4sLJpbG08Zb7RnUw3Oywo6Fc5gBIQiGCk9nWImj0K58Th+ec
KJ23GIwpT+oySLnW57QOp9di1D+QQ7iYArhxn4U6uEJYgipl3NHiMu2kuVisv5HUV6cKrOXElShG
UnLkKdXJAMZwuIP2JDcLPmebnp1TFOiunNzlJoFweWKhmcCkOnlQ1uqdE2AZ9V3UVzgkGZZTGO6g
tCnfm6Xle2nEBaEP8ChW8zFtK0BD+FmI6fNBFfN2rTzsHKEiuTySbe1lQFGx5qzVz9MIQfKBzRDp
gRTT4W2W0C4M6fURKo2uYMmoSKVqKuHdcAZ47L5w0lT6VGS4IPSkuPRFfRJaDFgMIBWt9lasVA8y
C9SGWEQNvkHthFbXymuQsoI2+zbOW5SOQPGpRySgPWn2KyoJZJNW8ZvWfYvnsQvGCSxjI4W8RHH9
u8XbHgeDk+/GIsN4/XdYRpWu2PBth9APzTdfLoKqEsDMykdhHNB9wjGcUY5SCd0teibWJD7BDoJT
tCx9V29a3RZLkW5Se7+rBt5MrTVYNFx1g+tA4nmbkYWlgBas813mF0KrOeGY6Eu0Bz67ZXfJN/F3
n67N/vXbEeGYYI1Mz7Qwci6/9tI1DiXU7L8BCcUceRSOmzO3N9yZcXIPTvt9kTjr+V8TZHXZLr/v
aizF4wLvb7d0dYCKldKFjyJKai5WZ8xytzXrHVM3QQQ3iL0UdYUI7e4BADolD5xHSJvR8Znclu7s
7xN8sy+k3shkacCjogItELy0LHbJwFAnr3Gt+DFiLmuU/zOVEToovj+HYljW51hX1zf9wCkHqX55
lAk3cAwppNuW44RDkkEgbhpEl5C01VLBrCnWsi/Zt4bWRh3HfMzF4IIeH99hIUhLW0NouXgh3Rnw
51rTf7dBRAaUZYWz66ltALHCC2tudSFO/nlOjvu4wsY7u8Rimo/sVvEAOR0QkpYx8OqfqRY98mm0
sQ4lRqO/tMBuqIKYgaN/WkqNO6XA2XwBCPgrrzj3pYK8cTd7SrAHRm11ph7R12qoh2ZT0f/KFRFS
NB+kKkk1tigvrrUwbdfkfmszxxzZ7NUtONmaFlG60/3hq5nVTW/Tpk9mTyWAsQVl3RDrNus/Edtg
knnu0Z7nwt5mZnK4K+ZMXG5DwMR4GehAZMqt2oOGXUgF3Mrney/wJaF05mzs4/Y92eZUm6zASPwv
JUCqB5d1nJsEk+wFBrNpv6Y2RfBssq4AW/GYRxAPxq0NxGeCjG/qyNE/yYMkEon9kASpU2Zn0zn2
25+1Y7Cz3RCeSzinBNj8DzMEUKF48KgG5zSZTbK5b3fchZeGNIFkWr03fqh9d9cLyiAYJQcfndNu
hY2emHv3LUf/ErOxlfHypp0nrpFoWyXpG1CplgKl7AhNHgXGCh7a/TyomZWoSVLZEO/OoPdhTq0s
YUy/fS3SLZWTKVfbDfuDcPmfHrfImVtWEwcmNYvyJleiRHVitd8lNpSRe1Btgxfo/Rk5ElDY6LLj
/HFoxllEZWWj8LAywwcjzipZ1GiY/bpV8IEIC9n1QNPNK3srgM2KUEXRwW61bhtNwy6AYIlk66EL
q1c78Wm2c0qTeinHmSuX2kfjke+Cvyvma0ak1ZTBk8mP6l3SkuFKXzT37v2L2HXZDkyUQhwbfHq6
JwkSUYTNn+nmBblwdimVYzQIlUtAKUuw6oJbCBFdZP42G4mfTHkGuXLhQCnkUD3JfAQgRDLIMrjx
MSn0d6C4wK4MujCVEzdYjlvFdfIUsQjk94DNbbqTAZYJFW8WmarI+i2IfcyvskqHU81DkhxSysfI
Tn5sTHfrZJI4/ceugpIsAe9wdBLRCZAnxDcOtrGN8K7HWu05iSQw0HmqJk6c/+x9zruADJ7Vcvzy
BvCAwErLAJTwxcPCJ+7jW0im0Vhn8L5DZwEIphf1dF3NxwVyWTVWC1yz7LdEaEHXdZxeZUSBWIsW
M7wJgXaDS0rDD5M5Ep/G1ht990oq4q/x4Nb3SPM30QNW6bMiSaG/1wyVSQjGFbQGbnTBFPBVARhY
Q0oLMdf/6LE7zNIe+Tyy7FAO5+Kr7EicJS40jVPGmim2iq3uvhQnIAZN2rWZHg/p+s0OjrYmChC/
g1kSS62ffOcRk0oWxmDupeQildG5Y3zB1QAqz6v0UnOuPsSzDJ9NQUstbvGJ8aKng/IhzCKtnBfI
Ky4Z+P55UJ15+gpFM7XE6l75UPA75raoft4y90oWUIn20EB+dq3pg9dPf7nZxzrpcMPrH7bStUiz
Ra8+sjrXy0kpokTMkHo8p9LEBkYRh9Kg1zU6YpOO+zJHDnIiL3bouOOvXKvxILJgZg03qRf4voJ3
ToAsXPApzLFk+Kr16Coh8Oz/2r1pTfxvJWWS9Xk3/TUPGI7WrXj7x2Nbmod4C17/TlhlxvPV18Ze
fU7lCrUImjW45nKytu7k7Vowg1Hgh7u4+ZTBSq1rE0rQfxi0OyL3pEMt5i9LszIjQZH7V6Q+dBQB
uNNhUFTsm0VT6H2bLkxkELktUY5FTV9hsXYWDMvCt99YbqsIGUatxPhZ3lKQOoxMzntRlC8yzv9D
R0QuzMbONPDhMogYoO7gpWU02dgfI9LCGEoxIxkebl3ziLvlI9hgz7zCjajKB2d/UC4P1ROXgnMI
bPl9fAjl03CRWi++0f1fJvSGemr88b3hNafj0mO1JU3OEfFcKX2jS/+/HmPHewpjk9l5oi7aBYFO
dEs1sK8nsWKkEyrhrGiJZ8d4km5KdTAf1ufbn+m9rGmQgqnyRDNm3wBCsMZCnvcxvXdlZn/nIJ0W
nm3ewzoolnmDgV4JFrrEVTe6guEjSK1/8/MkPDbJGTQewrd4L1ZjXnLUpW5yP7rAobG6eilhPQDG
zTzzTWbIek/dVScxpmD0onzqQw9dAyzJtDjl2CdqGe4NjKCRvwwhFJ0WOSLf9dZRYb1lqYlHpqLg
mVLOF+lh+YIxBvR3UKwdfIBG00OLE25nwRVve46x2kFNAybgf0IDXQ2cYV0YU5GTNiCyndhBz+43
knat0USwrKis0Uy5LVIBbSV53nj+Atc9YY+nOo9cuSV2ign4ssd7lavmhHUNvCgQfidV4e+qZ3p9
UIEHax8u+lKa3vBh27G1G6g1qZ8af5K8hhPRWuBgNWarKT8iUoWdlMkAlQ8+9NJiDTEB7Kyni3dC
fAqQC/fswYAL0ix+Kbg+O02qbCdiddPlJ/CmUnJbxBiWKSBHZbjS4PIXsT4Ybj1VMnYWMVfC/FVg
YYbKmJFuD+lrfw5U5NEq1LjLg5N1ZW6eog1X8d94qHc1D9yvv261iwaV+KGSwWZmsMxSNXLivquM
p9LfoIvLFs7+8J+kt2uzbOf+HyyBd/DQKaWr/XhxIQhqZqphPr9X6GVEbbWF8Ci+gk5n+9Zl3gYk
LlrwX5gt9GA0Ob+cle/GKVLopChBWQOp7n5jOfY/JKwdDLhrjK0Lv/hTF0bdfxBFCgD60TJVBS1/
zDqQc1CYsvYiwjyXLYf0ufsoyVokmymrREW3nNpozT6yuHILC0/YhjXD3tEcfMnQymeyj8Hvqr1p
RC4+oTH7w/gnIN862C/xyYqOqwZBNv7eBVxmwISl4qQIOZtJw/6ISVzhWQ+K9ZjDFOMb4S7o+s7x
8CgdTgO2ts1r683nffH9oAjxvYdQkB933JnL3yTkPT08Z7ROx8mbtOR9neXO8KvbpxZz1xRdNI2G
l9RmEgy+jSYEuQvcdNpYVL3I3B3+b/N8ZWU1p9HRYY9SEii+s8cxggKhPBreqYVCt+u4a4rFXY7q
boQAZs+8pan8WfLtZOYAQkXKTrGeviigyRjIZ6mLrjPxrPOXfVaAgvKR6QshVD/Rag2sET9+BZQ8
UpQJkjhRXReOK4M4lw8+blYW/OC9UhCf+urn6ty6DPhGJb7BcS21wWqOLOKperNG5r0tv2yC11GR
/5rH+Ver/b6wx6eKy86NaGVXw4FAAjpwtUgs7kLVmeYA/PS+tdPhXqHgFrvVUsQsKGFIZ8koFUaB
aR2vxKQAY1S1cnqwX31zR9SwJBPUJlgkwVORiALXbVOvycxXNYJWb9+F3k9wAV2I+NVqorGzTYd0
5fJPZRStlnC9FPBRd0WOVuwKalSqX7VvV0HA7k9nCV9+wCobyjZLWJBasFOgUafVyo8fDwVcC7dI
F9gks2WUjRNnkJo3Bf0mPo+8qcl7372sJ9mEFYwF7ZrWYlp8BJXgeflnwdrbl7yq7X9zspF0jWI0
OUDugjwkaYZTV4hIPc5mZtRt57Yz+RV/OsD2FO+hbJFgbeU/FJ8NJ2DgOUc9THSb+t1jzayNMRop
bCmKZriVVc5TkqfVb/K2uM+lPuxco7DSPl3HUBXEheOZyTrnK0ICqPAlstw9jI+0oM7cv2WumE8g
BQ3yBx1INzsHJSvN/3SBrvie3CIPplzek6TKNJVr4wb0h6bnxLt2910MMx5ePk477trl5YGHVrDj
M1hnE3wQ1ocgL/wkUaZrq3ej0QYq66ShzdAceKpKhFSJOMGSvmt3XQ/PLapp6oXD+QMEEhguKWNF
kTDzfE+8mUICkwDfbJHZfUQJ8qHgaQi5Jop8sS7X93wkEWp9zOGhFVzLitBOv3+C50PPStD87YBg
5m+o7vLg0aPFzJ6/NELLO2Sg3HquwgDFfFs5yh4PD5YtaJWULyXdR0QZsFErghDHldCvYXV1f27c
KUM3CKROdJdoaG6FpGG+jDzz2tmS2ohu+ur0xskBoDnnEbnpkD2EtkbH66ImHvuFipBRZytsj0Ib
9PhhcQntL2z1eLbtxhZ647+1os2iDjYBTE7RZqdcxNmHwvO8wsSjEe0U5ULqiVdocxa6sfD8kFfQ
xMYzBrvMuwWXz++pUk2B+7aM7S3rzK1mWq0RMZUOC9vhjV0uvzGxS4vtJD2thrQpUlUrsJnWkG9m
7w/DKXMWMVJs7hW0vI5RyRLKHSYLvkX0xwdnEzSKAcwY27Pkm8md6ZsmpgGHyEisFcR7frYxSyEv
68phTajhGT5EA8JZCzzURajleU8RfySNDUtSFEAisr3oy2Y3YVsZZ5XOSkBYa/GGFlhRnsap8Glt
LOEoNwyj/EZ0gYrPE0jnOeTQOcQ2Yb32CWVEFA+5lqcnvDfWXgOrU5qP5x0APzzD6XdknJ454yYx
uWexOT5M1xjusIGsUNL0Zh6oyF1PcQThtG+zF5vTHPa32EUDJaeAzqR4dKjaju9m2P72dpVShSk5
g0CV0udI3KFsqbasMZ6FDr0lEWpFqETfP8gokOk4YU3nTxZuAO/nisF0jhJd4wpB4J4LkNiW2dF1
jW5QXE4JNtnxB233EMrx8MIq3IgRN/+J7jH3FsbxuIIymwSz5CNKlhAVmtMO3yDvyiZhwbdaXL6X
HIIKaw3h3Bb0NXWf+Vkq/thsY3XOEQsGqDnBClh9xw8adIW8fdFWniy0ECaOH7kkPs4UYZkCa+Qg
IT/EWsp9+bgsN881/utK5Iu5w4Q+42sF5d73VFTBLbmS3BLH8k+4c/LYgY1AkRvuh65CX3TDEGTp
0sESTEupIAmrqqLnX0gShPtpvRglc5rgpoq8+VHLmwpeqI+7hws2O9qBsJe/ZIWS/U6x7UNmJpBq
9ZPM1Jr13y2afNYcFyctdl4HyVPF+i2im5vNejWYp+twM2iHTfreyQrN8o5448daiDHaYI4QY6eJ
8vsB4wjLL1Ttri4tgBrpHmCvy7MdlOll7jhBYUB1BIOFCNlzKlUfrfEqE81IYXU+lKrP7MS8e0fs
LgQl8khkBH3F38mDOwdcW2T2LmuDwRQWxS+1e90sWBr27QKZPzSzaKka0gOx/QsFtemqRsAAb0qt
/XooqSdzKjr4WmizQQWLkq5ZTaLfMApYxXS8T3rCNumqkj0sWT25t09PkpuB6+L/roL3MSMXcahK
PXvkWVhdna4F2i1zqEHrrdIseGHJMa2JwUD07NsesBKHGsxxsW+jX/83OJmyjqgHqMPjdbIu8yib
h4q3MaGhLnotSxSgcnvqohe8T/R6gGmynpRTyaf4aLs3oTE7/LuZbvEZ5A8BDjdkDoNu3OjR36iG
XOV3De2+KwNE2fy9twCeH9CTN8iQfxJVl8ZTPuhSAwCBI5lbRjt35lVgBRTGyDh+jpe/PDPvvmi0
BBUphC0uZNVMW6yIEisDDqadIewrciTXsIGejkqAXm9PMBF0lisZAXPSBTtMg4ut2OzeQNFF6eK7
4n5XJjO+qsSraGTAYtXRnFM7V0tvbn2532egaeVgj+nYGRla1A+phZoRBiYC/1z9pOBVq6uHandk
+i0AdRm+FX5bUABMmi8721Li9cM2mv+HJ0+/OHVb/gLnn837ugwlRt696XXyTc37Yy9kHuxNbXNT
NsQQ0lMmqb7src0mhgtVNw8za9cgV3pUNuf0ykM6Jcscn0wjejQVSJbx7Pl8gzqe7NYpqAI7YG0K
GXV3Cb6Xy7iaijmxGen8Oxh0iKu4ecT/lRIPd9Cqk5Z+q4TGRL1DrajZ+JG+P7WMpGtqA+EkzdeF
hYq2Y9uIYqQIgfgVi4ziF5kN0gPlE/xG6RM4Tc0wV0EiEiJeK9scYEVutfq8dncsNDshmgs7gr5n
YZFMVjNrCjXGrDbsqfHjjEOBz7VWQ+a11JKYfu4K6TRe5/XSlInxP3GLylSGpAaGd4Kg8NGjMVwW
4096qiiWdR7IJ0zKR64qVSRkF1YsUkGTKFYze33mt82LtXmw+TQ8dietEUO1Bk1uqliqwXi4bjm4
ZcD0ElCBgmp2eVtov6vgWCD8V+VwjEwVKr+vgxcrU5QomCkxfzPAtL7Zy/2VA/KQxjdgfpA1SKMM
GmUc0MbsUtSDvJzORK185k50cPyvZ0maPsHj2pMNfjabhpjhrjxE9ZTI+qvkDddhSBq3EGRCRf4L
V8bfGPuw7wpvdgpt7RCPNzQ2Q9OiPDiE0jcrASfSzVKdx5NCAOPD3WlQ+deT0NTBOesmO1O1WEBp
L+UnZw25hP1lVJZ1LdE9Qv5x6pVN87P535ZfmR6oD6fAyWGJBqMQmJlC3OoTz2G4PZ8VR0HwdODz
qDrQaQ2UkTHc7VYpXkiDkwacyjLZPI85xQcUq/W+hMJ9QstY4UXKFzm6R/ruLeFxvgkGhDwXbWf/
lRRqJQ34JFZ7Nm2AxqccWdOcs60ynjMGU88iqJeup97o905JEvoR6tTbyXQc0lbLtheRO7i222yJ
Mc7FyadAqIiaDPMPeRM4W7pDVRgno5sDFBozaFnU/+CaxYnd7f3zEyDI8oFwgxE4bSgzrr1GJmpT
YaFHbVpjo18rah1FCRz17R47QRJbYVME/CBbY0LKTWdk1MG/YVOvWKCu53qyLN+KPqOytSKIF/rF
2Zu/XXgCc03i7mi401yFd9HbUDidvHvNB5CV1YIXcOuYwTkHNR/XEqiYqXNKKR9PjjM9gA6Z9Hal
M2Si4Ccst8t8/InD1ssPp2vHZCsGdchex9NCZiGnqMhmz/xXylHPiXxx8eC9bqNEcmJW3W9mPCvN
DmFrib14HL/3Vv6jMBYw5ucxSML7pxjSFpLG8TRmlN37wxEzpHbOQ7/zbM4BTHYcO5LG3hYyxclr
r658cHqn58kfabgMDw4l5Fjp8R/ygcT2Np3QQrdRxmXYdP8dUUiXlxdBH0vOgUx8kj1sJsvgUWiq
BODmsO7itxzbgEVsEXCAEsYUEJufKdCZuMFPDZi3/ubmiSfu2/qNkhRn4ScGB5TNK4VZDYVpNIal
Cbg9FgKpUEsULgv5rYXO/4ybO8MN0M+hrsfDbCsr2vf1sNZzVqlKK/lih/mD+Gkr+yNy3UCDQISq
bnuH8ibn/tSkzeW8N2CfCIdPhbfPKair64snhJG1ci4j8bZJI/s02IYpUoxLQi4nYNm+JpkzizJk
B/rvj36ox41D54/YVcEemV1umNvJPcg4nwJseYHqhVrcye6syDhnL6pqinRwUGpXAVpF7zriE/Ys
R4nqlO7qKhrgInbgVOh8Fi4zJtofTjhVxEiORUT3MVAyedtz885e2RqQ6Ep3YVKXwdEZQx/zZ/Im
DdDqb8+4wM9klQgLrO1iLV5YfPOBt/YNRVeOqP/8rZIWetsNF7VPYinOI3pvTLYPlnFs6k5kiZMK
P1u6eD/Hq2xpu3FQ4fYmrSOqfdJAdg+7G2ck8YIHqf/n7YBFyS0eNjAMqXGZf61DxToH3BWcQdJv
yeVdeUuGNM8GiYvm9Oo2qECQu2hw/kADwYoK8wrzEtFyiDhS/8bU6wJIxuwy+k63QiS9mAruACu0
83sSeYxLlhEPPu/llyuD1mZaGZSUJAsRJIMIKeBnpjsQE0XCMB7DUit2sQ9YWOtFi7ryER/gOEIs
4fFFr7k5qkSHK2nFCIZGPPzFkjfN0i+HrM3RkzTxDK3UWTkMpk9YGEch4vNgu0nGGNj6WO81dDrp
Rtf875goR5IqPYKDOSDUTzFq6HqWTJdHjseW2SIMATefRItTtOjhDIu1OZzBgL0PAhT1PT50uqMk
TrMg398hK7di2LA/wZ6A7iIxDkjhmBlVd2mSCIWrG7dvBbG9HrD5U5b1nkgOWT3SESgGbq3t6gPS
gu0EJgHU4Abki3r4B3BqJCQTroyCHvBoqShNgbPQKMJ0x2VTCtGBJ9FUkoXXZPznWCnpLF6ONuay
SsQbDBQM7FUJvpb/+3t+ySspBMAaU6riEbFewq9+zsPNMlx9CU0JxznJ3WK6a7/e5ybOjXRau4HY
EXijePfJFT3x94D3GvspKEfM6udZH6/fWL6CC9+Puy6FrRynvBLIVYEC53kAAGggR6PW7zEtfeAe
xz5aVuY0CYS5HW8+xjWcS3NjmwWmjl+VYow9gbCzC14IHLzuN9KUsHqoZlr6coJH6kAWbbyigAcF
63WvlRoC+cDxuXkVTILt6Vn80IkB6omkjTlSifbJ0S5fUAmAO70qYgXLCTXrqpOTtTkOOGY5MzXA
edLP+RM7c/1T7PfjYmy8nCzRzLIFCya5+w024gbNeJ5vgIAv8sQeGp3EYOsv5lLChRLx/fOhqOyZ
rM252511LT8pDU8yohDMe/UbjRc99sYAxRJLgh7O41vnHxtLjMYl3+b0HygGrQyEn2JAaXKZ8inN
vr1bDp5LkXFYFnJC7/SeECt5kdD56/7HXHgdU2RZh6tTdUQEYaYu9ecESTobrQsBRZ2gFvy6OAU/
krEfgUqUo4e80+U7ZoQo4SAFzmSlOopKojGav0JGbmJF0S+XIDtnpXOvzeKkGLxIFTaJnhee+VOO
WGh/TO9KZhi98iq5gqZjrWk+Ap/GUUJ7ZEg1PWZI/y71TDkKWRwQ4TSj5iYzkYi7MNMDqnv5odKO
RsWxazVoHm44wOdTQXEBVcg8a+QfQ931bhjil2U1xHh7NEFaU0aR1vY+Bv5LANlNyVuNU++9SbVU
fBYXX+FmRSJO68fr9g5J8puhvi5zSZXaIvK30Oez/KUw7frHh9WoErYhYM9sd9qSBtYCIk1rFWtN
jTIgUXGCEfe9+8wHJiPuSKYeYnRdJWpjBUN73nOtNsZTL00Y5X28jPRKVk7Y36oWW3IPTblfTmiR
0biJ+jKf2uInu+Wx7k640yU9tNflJfAXOAeUrMz5IgIKjZ9eUB+5M8xZZi4+vbWG9uBCRHUje0BP
iwRb9qwE55BLEsyRaYBT09n6qKFnM/wCaT4lCswDBC4shkjZOXmfiHonF9qKFmiXxUdh3HsyUXNc
jvToATxIyIeT9fH65o7Z/vN8+dwpY5AoCeVHX7mFOGG/YbS/SCamp1GDvp6EymFnAS9NAWibl9U2
v7Hbe6ewLMVtbdIlKPZC0woBDKEda68/ervctLtPJrw+qkbeHgAodzRNtw2QR89X3HEsJvMpI6si
oqBq04/aaW2klf+mxRtEnP71NYn9BabBjN50Uy2acWJIIqUUAAeYx+x35w5PQOREgaaT/4HLYRqC
+90XM7vVUAVlGwiuxxrO5wA3tGAtv+zzCDb0ZjygI+roTSzcYXDXXzVto7RYNnkG1yTXjDlWd4L3
LJ0FQIPUapaT9uceBKGHuxApO6oamNI1YuszKbYGPgYc+fMOEUlh2TRcWGnT9KuVvk8Dc9sTrG/x
q7JXUVbreFaYY8Dk9XpLBwZVdCfTvjczhhfFigDuRwIduSa+62tBbe5+B0IvRD1qtBZ1n6eSg79x
rLlU6tgL77CYIEMIGkls63DTuU8UXjsAmrO0TkdZGhYgKFAgW5PEh56vC90QCAWY1/CDLlRUoxIS
kzrD+dmvMZsVGBGaFQBZRnckXC1aYphYNNJY+5Tdp255yoej6BdkUF1PApH+n5cG7uUTzGhREify
lmVhJs98yXmKiExvHTmfcuzfhphPRmC77ffJSamLR+yH4KQZfLAgNk5/CqgraH2bsTpEkTj2fzUk
pZn4qaZv6zuYauxvk3VlzOW5Tcx0keSKQz/swfMiXCz8/Z9N2vNqdewDq/z5FduJpnISo+GhU5w4
3LSi/1HziCaj+qr0XFz8Dqi/XYp2Fxh0i3mEut4JEHWVg7o599aj92QZJaulBQGiAxEjdpKvQIqR
0N8e27I7onYWr1zfsoUilTergNBNidUHc3+ZAKcuEr6Gm1fM+Gav6FoM33MZF9e7h6vhCnkczP3Z
sFJCDyvPBTzG63hEbY+Arur1MhQYs4pPxt6I6lDj89Z95ayFs065BFnoMfdgsZK1szBzFPnFGJst
xGqZ6ZX+CwSBUkFFhUF+XdWS3CELhjlRrCL5jBNAZGDSgXyI0GLFoZJRQ0BqKRC/tO+g69stJvyq
lIIcs0yE2hNgwMkAvfMLcV+kw+2lfEinWOzQnrGk3TZs8vdmETDhk65zHJ660iEnW7aEP1PtWWK6
qQCwD2LLL8FAOocg0bVvkdEvdJfAAfsVO4KKEsoVvOkDXG0PovA3JzqR2Tl5mPfX2Oe4e97svwu4
Mt5UWhw+3W/R6nGhi4lxaX9ogiBmhTXnx3aGj9UojZXucygw11ghLdRJtlCZ4WfHCcC8cQXBKNUd
SU4iuOt7+FL6FTp7qS7r8t94yizSlCmUGJKLXUWbpkFnPUtjZ+nysFZzowXQraQHQGdoMiWm8EtD
FlOGDkTIyFuZ/9ssPFZ3EUdT7I1FU+2fEX90zc3dkyNcYIy5VJmKpyx1Doz0IeMz2BcH+kPduIY8
8ZdpNF3zgU5qVgN0GM9me+nifMdN5dlpPtcbYuCBkPZS90NN5ILQbUQGFxhXQvzKT603CcW401Th
RgOEMkpEgc/5fYYvVC0sSlOI8t/Kmbj+03L4EFxEOloqSbuW4AVOp5WtvniEjNc+CqgWP9hYyZbE
1BjQXQK0Get/1jNKMZ5R6fvrmGxP86TaeaSyepaKrzEZi1djkdjyS4k2OX7Ad6P34PSs0odDNwbQ
BfEjmfNVEJJX03pPuDWOQRn0LwhkNYXbUr2GP+EbMTLLEbVPGqs6uVZQr8Myj2tuKhrp9R5kmW25
llbF30qUt+1KTlK1bXDVcebH107mK/rAqFFOckEOj3sbza8xc76q2w9ICqA8yOgTC3hVtXwIXThE
ap+bSIpRrYjKvZrd8OmouJVsOcBN4ZgUNXf4jqO6ry8GDp7N9MQsi+8zDmMUthBVz3/Y4w0UsrXY
rt7iRplJHudlnhjtacV6zKHWny2h1+FA1xe/HXN6RwY0WDN/Hmmi9vA+mUxmRcgcEi9Uq0m/nKxL
b3rUtjOtuNu0zQkG3K8o54UweL5il8ABUnDQagKnYccbkZ1t3FejsMj2tm2TqQJmr8AyXBLs54+p
VxKNko29Q3annNuk9huUHNYJbRtonzlJPwQuJ7Wp4FXzD6Kv5JfgukpgJovcVlYxerIhkritBr5H
bAbRwhRLvarq98UcgWMeMk9FFdE/+RajyyQMam+mRaQ1ftRZ7OBimabLhyllXgqpkGV3fqyQzhMG
3tfcJen+pw/kRdVHU5rQTFGTTIHJ7Pp+YDcMjIKGBGDI9+sCWGPromX1PDFVZnccRJ2mawG2wsNZ
VfSg02WzxEHEMwyW0BQ59k9t3Dve02Z/1EeyR3tv4e533m5Pvg9bKyWVxwkZH2BMpgdq16+N5AxA
PTy6hJ7ZtTzXR5l8D6n/gkBOwYaud+XkwIBnkReiF7qkOp3+cNw3AAoGNZmnTWuoE28h5Uq6ZnHJ
qXn2hG10ehVZ0/hzLl+KPgCK26IbPuxvazfO+ZtbvS7npvfw3ZcX9skL5ZGkKxL9tIISfBdh0adn
McCOVQorj3MGPUM/CIBF/cqZk+f3YNCArYSSrAUnxGuTZuzzUaj2i9itX153NOaylzqiN5pweoOt
k55KttzR12owMhy6j54KLJbrWlKaVIEHwB1/0fpLoiEiTjlIg0v5lofyFyZTFg7YKS2xwT887TRp
urFG+PfMSHH+ZAaiRp9ToO/VuFxQm4Cp+vfzlwHEfjJB9ua22lSscnRmk71SZVLe63KM4ycRlt2W
8WXdpgGjlS6CqAgXBn3gKMHtFrn1lUYgf50I6wq8sx5r98ufNglaaNCDetY6iGNlJaBNo6Y6DYjo
aU0fu6w4+To4ErYIdbEGAqHwM9BwLEqWYCVkmHpoMtrbyu2vFpbPZlCAjrncIHpvarpiS8Gaz/pR
m+ErhlM9IazVc9EjxFFIFS1hGwAwNMBj/G8BoYQPoYNxBzo/mwZIy160IZAz3PWFRc867fhr1kZU
aIH7PX6+8UY6kEk3d/oFxOm+AUV6toE0xQ9G+pu/gI6tB+/iIRAjuAEFvcA4EIGhmT6qy2ivlLVo
wD8IT/HxmbNRSZ4m+fKe5FEb3R5TKpxz3l/qbm0dESuX8Y0EJ9j9LeYxYwmA4DsfnDanVJo2XcFS
M6jqrW/5zJw+ND7oe73zuRSjSKyxN8pJJ7PZuWQDbLVq3B1nCY7MzY0FKpzuiWQFY2wr2OzKa9OX
qp+1zDv49mrsv0gt6Y2Rf/wrBM6+LWUcOE4WRbJwKbrRVsvxuajzLq83/b5sN23fKeJko+1u+gGy
XzfSrYN2lzIDAc2XxANJsuwxcItE2K8GVWojouLdWXTRXX6ZXZrOOUG1kLMvYLTlcxI7Z0MTyvI8
4DIJ8cleTZUs/byD6DhqXTOz0GvrXuaFYaJ+Yg24Z/WrOXh8x503D7byuU0i+j2lukocjd65VNWf
rGw7cGe4+6yU3Juq6joYVdtR0HikCViHeHLik/+kevueSur7SCABc6/SbA9ZwGuPo3rVg3poi1SA
ab9sxTZxFNNWSOBRL0ALmo7RyKPHdouEqp8g1sF8lYBwhqOkOT+6oeVrVMnk7wPB7Qpu3r7zeY2Y
MrKx+BYiiCW096KDUhIKXaNa6OWiDWeqSR54vPqR3O2w+qusY1tZD77I4EyZNTnQVBW35cR5MZUa
PZYXhVYUh+F9KMAP0RUi+0sAe0bQxbYBjJ9bhOikLMW2jvYIS2D0p9DVC7zgEuT4r/q4x7+QUKaE
AGfXDykfwsdHAtBP+gQo9ISGucqZgsiWAP7jkQ3mQRPdsY/wA568T0KVdF/orZMg4RuzlO4JVBRm
CtyR7+nkmcaiC7DwfFquAZfa6R8H0nNeNq/exilLaNV4wHtXJ07rU0ckKbyXl/zzPg12ydZhhI73
GZnU+BP5Z80PwJPJ8f/h9q46HLnZFp0NHMjtBqyD8uV1Cq9v8nv3yJdGq5FBODNvt5p4bFTr/8WO
qkcm8ksnFGW4MnCt6m7+xc1rISFMO+ZW6bLYlCauQYTnBmMhiv/YaEQxg5DGj6gT4TEjjuS0nHpR
2x2h25vfBHoCQ+tAiTbYnXjJz9Jbjs7Erbus31hyAADML6ipgHS3WU+hXnDKNGHp9458WKBHYXsB
Evy4wRB1ErD8vrEM4VsrIJ279VQMKrS5MY67Hgk98yTgbw45p3phdP2586AV2JU8LgDgZkce5jW0
XW0cMJMugmO0lXNzTMhOeV/LuB7DD/FIzGVR24NFlFCvuMggh+VuqLDpo8knweGbwbiJhUFPqCLr
OmJ+R4FmNtEN/ggHZeVCcHjmGGhY6+sDcDKdTtI6N3f/gWWO1k8JNnqSR6NC1RDbg1tgKb34IOeF
MIaySXhSkxKYkpumUpYmxnDTGhcUNm9lzlD2iqINd/XhrAhy5ZCEDFJJonBEg6OhheMOO6+oW4wF
Zu1TBGOKXoTHCTDRfdat+O0oVXmP9+Cy7efJ/9UcrPTBCwcW4LiNhcfNGIfRtBb+qI9CQ85tpfyS
QiKIMGVVwMcPyK5sxyjvW50P/UagVxOTnO4waIjIGfkqHZ1XhPqpoeN7drhT44UkqplUhRkLT+Iz
FPjuLAZ2tqLFo8fa2v8dc2zMveCreGrA13+7Es393tVZbAS1KI5rrsaMh8S9RtVm/DuzBQ1rgNTK
z+E7gun4q1wSVOJA/lCD1BQgP45dicwy/fcd/lX1PhdlqPm0PtcJZTWZ96S03zrMmZF3QNKXR8dt
gQ4ZrRYbcCqupyoxESNE+kjhJFY98yBu3XyAxnXLWN7vJM0Nyl+Xx9s+w4RpAexwdGIpUdTauwp/
tEVNqaP+akXmS4x7OLI8D8fatx+3VfdGAn/oYq/NvgcpyDvCW5jUYGlIvF1ge3VtgSxRQDcNXrGN
0DUb3FjbYRSj7L+wQEIsRRqPj9eld/QeCOEUDDqtUeG3qghCJBujnsCsaR8qBkj6HuUMWxpOpNms
VaGGKCItcmbGHDjmCuHaVOgcCeOjLsxJYoUZ79s9aXTodLpfxIh3LUFMYLoalyutdrPfM65fhVvY
z0f/f2+A3Q6y6Vfyq8kvMP/w/ulCHqL2iAjxOnj7okF9Rk9A6ZJPD4zBX6VSqSIJwdC9MVcCJLcF
mPOlgQ2mXtmj4AD7UfL88t35kX2AW/zyTWFB4sWgJGIXCAnnYLIoBZfK9cjkt8+WwreLXRVcVvTM
PUQkFw0WBQY8G1fa5m/BLY73fGrp5iK0dZR6170GSM7ThRpyRWg75NL+IM70+KG2aSZ+pcddrazg
Q5R7PX1el1qWeJHXNJ03F80Hbl3JfinYt5BjkPAUlXaeg/5vLMH1SFTm7u8lhQiY1lzYpngLf+er
wQNDupT9m7yxu1kldNiAutnOgr010g5iPXxf5Jl4qLdVoPp339xzuyCyay0YTYuY4wPTBIQkNjI4
AHZ+5Nv9XSY20NDIUs7vkZqS2Mxz5ZppxeqOhamUn7zBUXplSJ5L2ZV9z58xJoUTHFl6E3bjZ4RO
VfaZljLhud/+GZlW1f5f8q6RjQ/8N4GgjkxihkIJguLc51tqNSOhYi1/bypk3Xf0rb8HGD9WYMvf
7NMHADrdFYWdSpx3OIhys9KVo3zR/6NkMkyY7K25OlHlhGnHQeWF0RKz82JciDBf2EEYJ7fQ3q08
QbVlw4lNhXYtqAp5CrpqDInTlxxBBYlB2n69u3TL/NfZnYfTR3Qw6XBSCVNnFpU9rlwraj2RK7n5
MrLXdXjauo5QB1STZNuIVd08kg7k3AWK+KIfl3ZS8eTc36J/DZfsk8MMluq+zYV29hE5vNPGYXqv
njZASBA1ildVjS3TNtOiA4/l0ffRhly//pfKqi6Kid7tpM5hA0rnRG7r2BT81Z8CTAXTh5Rc5cDb
m7HvZNRC5IfbvKIyIMt/sHKZCaspFFdauYISWz3ovlDImlrdVzexhKw8aNoHce8Kbp1auF2galrM
RTFPaq/BZFpqbDyaQ3XFyqGkqQYpn8HDDuaJhvxl+2N00kwm5AcJGKLdTLRC6mtnQKV+Id7pXRrd
Il2yFkxKhc28QAjv0XXLWvR1s92nSI4fquyVARzDgAAwqq+ApFwFwjk7eI66hbz4eeLVWyuCyjf1
4KsBrPIXMgYcjwbzx2ucr63DP4cib2OkJLBkbUAwJ8No+ySdCSDoPvrp2Ymay6nSsgWfFdiPagTC
m5wxVYzDWGICH0iIV8LN7OWcnqGwMl2IuFVpbpCZI9h5aXx7M763xeJdrtsGk8/KjyHrBsA06iYT
0FCmTr42mFSTERz1uJpyK+o1cDiH/zqctgTHbRAJAZ+s8kaKACV96IaSTll5qFLP1RhGSGV8ies+
JFRflLBbF6sVZQ5Mvb2jZd+LL5lpYkdQ1+S1ZWXEJUCHbQhwEAAziEJiLdQ3F9l/QpmvHUK+3noi
u5sqc3MbpwzfO1bRwqGUk8TlGZW1E/b9pQ8GnrZKwhXrmIjaYHvUDc3qgOl9iNNkD7FpDlWSzl0c
QkH55mB0bg39W0GCGfltGHBmMiTTv6nJV6yPgF+jjoSeJuUouwozeQNbIzD2pjMQNTW6ymnZGBwL
oSbmBuNPXOQjXCC+ALr+ZmsxIZGcTREhwcHeqpR457npAgleb/7bdE8kqIXGNaDj9hY+2heyqZCR
Po5RMR8cNcLgYViRm4RzsrfVDIW7F7OV6zIZ5RbzR7ZeeFhBE/EiA3AdGMZNv5PiI5Et2kkwpDlP
zmPt6Ekmezwjn28Deh0cHgmYBmjKCWVjT3+Q+CZImtelYrifHrFXK7rYy/uMkxgJbPRxS5zwEbNW
04gY7QMwCc6evtbbqhIXWjE++5EFWHiClq32UpX8D65i+EzOZzSIsVIRvAe6GKSySev73FVhDolU
59CA1L8UQDJL6jKPeC503fQGzlSxBuV9XnrFtESviBy+U0APjZPJttCR9nJik1ie6nNqiPIsPOia
0xSti+f3Hmh+pRthUpVT88wNI+hwB8XNpguN2So8EVgaRurO1Mo0XqY/XoxaSDj3GESQgQPYqkO/
yjGR5EQvVbDD1RenzOSG5niQpf4AzVnAYr1VTAEsB8YEpBpyveiMeoQgCQi5S15NRzmirzb7e5ze
Q2leIHULsHJb5b6RhJPEL1QMXeVEinopH4VZXdaNWQ8VEgsXxwEcLEO7gBO08nJmy0lbrOyELPAF
jYwbhKpXXZHljL7HPR+rBD9qm70JiTX9Cl3ivroQkcptCv1ICotoe6NQniYX3k0/o2Jh/BOtGjWE
v0oE06Qz3E65ESIVIbBWVCHkNShKB9fJMrSaCZdG4JB45+OZd+JPjYNzq3eh2EK79PpiRAByb5Ns
yTxzoso5HgNYWVaDkmGzSycp+pr4dMb5GGJh3tWrhbiab7MXRD89WMUW0apInG1sL5dLFOpVcXVo
eLVLe3LpxaC752bsLyngqsAie6lfJrLHpylKwNFS8kBCWng+4H9nCi5re011g/hnKYf0uVydqGBb
Fcs1sL0GwhN13zgMokGjinuQXl3MoG1i1CgYOIYuliCJF6YWiLxQ5Y2f8XDIvweYj7pXuyuvR+kG
7ghytVJAucoJjcIxOFyYehXnZGC0PMEiY+u+BGVF6NtSq04QrPa4vDjngJ1IK4EeT1lSgGV+gycW
D/U+MCHYbeTkpD42ZQZK4+4fszUXRO7qSdWEaCdqgEUV/0T3gR/hhuRKtO/5GESfIUAbmfR278Ut
5tonY7Ca2GrCBqHk6psjKVwaLJkk1YzYLRlH3/+GFLmXnwy7Yp+W6Uy3GcFBJUNB9VKy1Svp/vlW
45YRl52UBNo7EklEgltxyacBZlVU7D/cIFtIdplc2PWvA5xB7dFO5E55WvEgCDxUPUyGYMmyn/Qx
cErydZSZotngNlaYDDx8VGHrV+THhG75u4AhlkDA7/yn1SM56uVi/RfnAX5L7BXaWuSxmdwU+U2o
HZeRGcN+mAZJuGmRKL8rOFFwXjE/Hs7HJHREWaoDr4PijdLBovnW4ORRhN+TpQDv0Vb1mwXdXCss
4ZLuDQLaLXGuJhx2CTdy6Ut7UKCU+oqo97jpHFhv+E0kE9S0mQekBdnqJxWCUe6j9vYDXmfEusds
XNb1O8bDM6jnAfh2r0j092gSvB0mJPFRfeMW5R1qosn+3m/yASKnvyRBWvarkUT5Edc88+P33Di0
vbIgZblAa82BvfpObbPUWvkswyF2FQLdMFl1Nq+OL59ufr+is5cbtyY5b/8GHpIH2vPeY3rzyrbx
Fizei3FOZL0GeMEiGotYJdao1nHg0p3lMajpWWxdO6MaAUvOpPyaw41fTstS5kMekJskFYgLVrRr
gV90tTyntlAYeSiNNPbktJqST/7zuJGXVMcT1XUTvtcrEoRpbx3f/i9NieL7RFP11NyH0Tz8L0+d
5uDbXr+nZx27mX3nuT8WkXh3XdSCiIPGWOGaJvx7J3+vva3iYsiAYnhGKc+Y+6RULpZ6qKfbfpyt
gIAvVuV8mB+FCtcM9/NSJlqBS8UfqUbBoZEj7CKUX1cP125yvWPyf3BdirDRh7xaVo02GQf9VlhH
SMZNLdhM4uBKh7sqDaRKt3s5+qhkCLQUTnEgbhdIQfPVDvNTCtWe9yosjV6+BKf/DY3SodjZVjVz
6z6NBqlVR65RL8s2OJvRQUhUKmPmconJO/XcI1ZqlZYI32eNerWz7VdMWtemqhuWdX16nZJ+X8Gt
gxtdaok8vwn+xNC0Z+U/cUU3T2OjUjMbdWuL0R2fS0arpCfqbXfr1C6jKrYZ9b46NKsPfSy+Tz9X
j88IPdw6VXln9yk7IzEz35C1kbAcJi0KsIuFOVeuhsZEKak01rNBB+f8Xi9DbwaK24kTqlT2jdVV
CBr8zhzX2+SulHs/IVNFpDTchNsRaGLgfU0NkKs7+auWuDkbDMPEZryGQFtKCqJemgXRczxCSe4L
wIAdx3l2JvGatgDI0tzFpUFYUGsZ0/OOoc379BwvCfruSDt7lqVU2TKyE4cSJSRJu7k/bz6hJdBG
DQfuYpUETHw0HEvwJ8XyyVMdqZt8YLq4laesMlaiPn+u8BfspWV8oIUWAwtKO6CduFepqjwV706q
OxSTUXbzXukswvwi6E5pkrVhUWjckUm9k8Ff16mEHFWv4L+Q3+eoUuSPzwF+IzFxmIzf7Bd4uSSE
RGME9EbV8PX9USpJIm5xNIA2ZyfZqRxh7UOCYJlRsVs1biSzlqYS56e31HCZCvnB0sTcCqqq8BTF
3nEDePcPdZqwkzEtTwP1tidi/oYdkc2l/rEyDLbZHI7aqlhkpQ6EWTe6I/HPU1E8BpvnL7ue6Vkm
g+jSIALXMWJ6YcdSCR998kkIW+gPhtUr5ISLZozjBCaM8XyaDM0bDYECNkiZgrW0Pa4UddBIrH9l
mx37/scHbV0Z5sXMUl8K6u5IJ05IFqDlWc+mYVK0pH7L1atQvP/+Hh3nWT9lMDyYMrfmLu9LnGJc
3MV3+zyKVitc350ktxKrKRtm/vmBIDStKOLDtfZaz9Egpf5OUsNjADasf5kM398v30Vh7TwWSe+v
iBIkZw+fjkMzTk/tOmn56oBHd4ajf6huGzgIxNWJzb59o6S/9IxCQsQCN8RalfPoiYJcXCWFsBiE
hPyqMoXEN5jlQk6RDaMtwPOkHlIFf5mFLeGkMw/PQEAGJrsnDxUVHwoi9iU2qTSeqd1KvS/NfV0h
4m/ilc9kgMvWTgSlhB+0+uI8IjsgOHUrIE4uBPO2F3ooow9NY6XJ5cTnFiJbae9DYkczW8bCqz7z
+/FAVKAkdsvlGJeC9E45/87QS0r7FMcMbbjEWa2HuODJoP/1Xaoo+nB1/J0W9Yg5o1FIbhBZ2VOj
fiH1Bjn3qDDuagRq0cHmhOra/B6AxzyHBUXZDY0NusN1NTCCpoFTrkvfvbn+0z67zXBnjNEqEXfa
/xke+waRCmKaBT/wPYejjKaKMDaL/3yo9hKGVrXNq0RMPnfZ+jX0sBDU6LE+e36X32XQgdnljYOv
E5BVbL7L40rcyArlHhUpBhGPjI7ub3d1nTs0E3yeJpI7wQkpsb+OKze2qzY/0vIlFs1DhVx9XzVw
QjQzcQIC/Mhp26Dxl5ihJ043LJLBnERzm8/CvfQbL86gHIET1Q/RlkhqvAWRPtP2M+maHtqHrK8T
xulAmhxtBsO2pvBjRB8K45b7JdAfvJAckfgtjMO8QFwPxkAY4WEoqTchJeAzoXcGiK7T+dOPqYgA
MY+bWfMoO4S642ZHsHv+nhH7dSyZHuaDTfsnjcz26P94ApLc6OFIoUyfd+uZSZCM7AcVBh9n3gCA
C2Yy7TVH3Na7K+OGRsqF829MV+bXiKCJt0l7GnM6SbYnnOsmIblu5rkeNcVhUaI1HkZcWyB0ge8U
p76qczK1Bt097YUzFboVGwiOdiGesoTNaQmtD4Z57I7axF7iHJvzC6ce6sVdVK2twEUglTILGND0
jHR6pOLw4Ra3HC+DrGeyabOUcbbjfnfmV61/NRlp1UB0AHr1cth+ZUJpjb91K7SBAlAHoZsLO0r/
BEvYvu4VGT0R2Qo9Fyvm7DRy82GieHA6Odj6M9Cyms/d3ZvneHaOvUW9xS68+KIs0goaEgM9cWvJ
QvE+3Vy1Ouq/P4mxZmBfVVZoFREiZzr/c1+SlyQ/gE3yZC1zVzvsp5SfZ84QSs0EJYZmmljUSAPS
XYVxmk6+GTpj/q+xT8gUVdzkYxTOlCDMlbAW9l8jS6jGUe9duxoLFuUgh0kBJS1dy3314BY/0vVt
v4KfescqGP6Ug6UkxMiXoPX1M9L0+k/EeZhyK1ys43oUiq9Xs2csT/Bd2s74LApBIwCR3tmyYJWt
QcXpWXgg3iJtNtFZWWy8Q6bK2hfB6mGmkwKvVMH9P3TaA2xmqkmADCNmI3X4KcYaFjesZGkpkEcB
TeojOj158xmfBjQMXZS0es42j0t6HiReOYzA3vvCyP3pm8aLBjPRWtOhmJ82H56SKVYxu32KerDJ
/TLjCJB8wMC1h620muqwRtrlxxeXnoPtjFyGdPp3WEYcvxyHsYgpOUMeI4Uu9oECFqB9nEjoh2F/
Q5oQ2qJcR6Yv6KsxqIpcnlT5ia4oW6MbyJyzPOJYKAqufcyQV9/tx7G7nECh+ycOaYXMPAioM8jd
uy+L9DpWj/PKm5rnwDTN4sXHkmmeX34S1Vap2ayQhm3oOK8YPcf9094yztcGIuN53thiy2WL7nMG
RxcIeRprsd7Gzeqmpa8fsbPRXSXT/lnFrC/feORvlb1F+N4JdEG2QMoSi5p1tf9iLRd3JZdkBnmV
iL/Z4HCP3OYxoxUtaWTjXQ6iYKSl4xp+i4GJ+BbVnFgkfqLClFQF0Jpgg5te4DzasnoJAYvmE0g0
lc2J7EHPGjg5I5U8GUtHIbxe/1MDSSFQyZziI0YUEvuSGCf/4GbZSSR8k3+JEP4YpnxbvAHNYFcf
yKFLs3/C9iEIWLgVK8OZQvPD3hKN0dssYx1V+6pD2dY8k31pgjOWXcJMdmM7ZRlaCRKmnSE5dcxI
8w6QHepHxMfgk/H6uipHcpWvTFjb0sN1MhfsWoMHiG2+tiSJOYg5Rkx2ueXQH0CFD2w1Bc232GsR
wvCI1jm79sav1WYoMlLORbalcpMbdBA2g6IdYRKJ7gN4rWAIaZ9nlg0lMcFPiJ1PlA5dgnHJzgPG
gcZMSoWd3nb7W0P558/zUu27oDsG0+YlqTxQaQUYw59sByKZ7ioVIKah72Z+uuVI+1e5moBtIj17
SoQuWNnyeOoDq4hhDINRMI4f1ywsaVYiKoeiYIAVBCHCRDDsAalpVABJF3NhvVgVQapX6yhpNN7T
VFS17Qx6xNahKRnXoGVwh5EvN6N+r8OyDoE5qzeGLcUKiXKuW1pGobH+HbZv+5+MEFsntawuRyHo
S+cJtkXKJJRU8sFJbJPgHhDvtgL4KQyiIvlBmDtL8+GDxKR5xK4uSgMy7P4gJQMDAswYsRb7ODUI
T2qN7xqrQjAVZh8pwClcfs1mUtwpQUjSNW16NCzAWuPKqmpfRW8p64Tr2qGu6iiw239EZ7U6pyIv
VCbV8qNppd74l7SwYktYQxpthP2IY5YT53dXMTpM2J/H23oSKhaBu3RskAbqFUFJWGmslaA/ToBx
d5+tN2c2hD8qz6popEgCR6LfieL5P7FJmMtBu1PAut03qQnwEaVNhepqgTkhR3VBMScliD3eyCch
vx76iNjYyShzHt4RPSjy6CefSu0+K2iOZhiKpz6DLTo3HDLxdktHyvfP4SG4TJNw27xlCR7BzKlh
ZUjMWVdaVmG+I7L2PPb6WV0f2lFmJqsvYm47zV0vhfVRlGGWzWC0J+t1l2f+pnExa70coZuPSfh3
Pgs3uXjroRgCMpOnz0eGLXZBLklFKQeXd7A+mI0DHp41Hwdgx04pFoajXUfMjmbNSMf40Iq8SOMj
pIz01Gd0CyL9iyoQq0Qx7Uh6Y1AZoJ2vvc/PXEZ5cb8NMxpAQUc3Xq3UEfkZ1Bm24wFAm5jfu1L1
D5ZBGDo5gJPcqbxPL2jwcCW9AU17pltdNznW41+PFP24uSht6qLBV3P8leToE3gCBVNvL3BI6M7G
o4Toxfj69H/xg0O/XEN1Ssjn4O90/M4wPzIXhZ+omSIlG/KOBoPH9K9wyl28ciJcMTaDoRV3tinK
7ZoWpkBF5c/D8XJOUucSjGW/h9O7jsnvFevixQVcO0+QphE/FuIAs0wsMw8B7Dh5bmwHF1sABs47
NumDSWtL9PSv/qPINVjO5b49W34jr4cANINxXKCu5JEQeQMfagOZG6V5pQMIqWUK7H1N5JmQwAo6
lcMnfrmDFLAq/u+cEK90NiajAaXO9bnaI+u8hpvg/F1bF7jRCw/J+glHh/cfPx6ACDZwyOmFIG9x
HNpcFsu/ysT9B7X+FKhMzvLAcY4kIDNKONC/817N/T2hkyRTZwsnNpV+c87WPbJq5uExs4Wpv4AG
F1uA11iPgkfLVQvOZR5k6GTLog+LyT+dYvA4TL0B+7ovEmvWauYDAExd4bIpPU2pj/18fflb4UlH
GMl4WICopVbCA0BVInqioZThVBuD6AQNff+bUxS65XcgCSjY/a+UPwS8WQf9LKYIJ4AFxCD80zD1
xiiMUWVCv/8k2ZJLStXSdV0WotkELRbT/CFYTv8/Zv4VihHMyMo0wqU13wKbZsqTKgOYXNCoG1vR
Xpt7SeHfH2g4wgEy0OhUB8vk8rFcrdyvIB85Bm++k9HtHOn0wUswqJOCb6EpArMfotGoB/MOUgfs
e7siRdimN8KjT/9f55iaBJI/p4y7bXdscvYOzNprxF01I6pdwcYuOGvjjqb7UnlZXU+UvZDHk+NQ
tWEWl4LB8JPwWQbgpXCbJCXpMbziJ/66jF9bXDSyop40r2p2b09deS4kzhCmlYXKTnu+LCjiQJRF
dav1SuLw0flqRLnTIe4a2CaTKL7I+adkfMry9Fwov337fB6nsSrSjp8+Bjbw0djrbyfsQlSRxH3X
IUVEg/+7A1bHTKqQTmeRWtiNaQ9R7Mb76hB9KS2XYdbPPuHFy+EYx0EVdbITe3/cjb8RTscQFA1+
nqXhBLmix7ep6vV64TiD7fwdba2w20o5ltFmDRQhJ+oxi9hGCvz4y5INBb7xH+MOYYt6DX8ZY7Jf
YQcZJ3N9c1fWsQY+t0878fop76R0CdcGCfcKS06msxQy0k4/ATzeRSEZGFD29xXPKB+QAVyGvmys
o/yT3YSqZ7VYzppwneK+GouLRaR4ZPpHsGM2BnWmcfw/vI+2dWERrK0QkJwF7AaA7uEjsINappAk
52wrU61AzF0pmuAhYZ7gythnBrhP4+D+ugUV1miUKyxc6XWoQVSZ59YR/g9v7x1OHzJ7cTNRO4kJ
OL1N1+s1rsy9KzJAyzaZfWRC/BaLofgCKSZcH4+Rw6ZKih/C8HETn8QpqBU/90dIiLjZMY5fdu+y
T870GqZN0cGe5B6T0gYdVga9vQQ7ZT+r97sCn6W8Gum4P9JxuCaZPl4fVc6TdFb19D3LpD2bfnqu
i6Ke8VzDOP6J4ME7keG8bMCvAK4wvggokjYbDQTJhmzDaetK9Lkif8DSpoh9zkSHxrozfzdKvskl
yq+4xp/pb9s0UYkKrMRyXb5P5cAaNIRmO7Pl0cPDHg6v/FgglI/VtPoUN12UC9eqqCG2lC/SvRo8
ymq3SM7plnlNvgfwJ1gEGc4GhwXlzygVyjQbU5TOQv8skQQABuNQfraeazA3N+x2A8LBqq6OVxlO
g1+6h6PVq5nan1E48yE7PgPwVAGUi8Cyprst4L1P3Nq7dkVRu9ymZrKMkCoeOem1/nuaHQHj47AV
jrQXH8jt7ZtaaoVm0mWLHMxJuVi+KO28S7GO5KFZovnpLr6t04ryJSC0xImFIHkGVAIL2YbfmeJj
3XKX+cp7kuRJ5vPmrFoHO1dvssWelnAM3hdsHPQJI/VexDI6nid3BeL4lVvaEyc/YKGLusid4DY7
1qSG+9F74scaTzS0M6upQ4ntNyi4ORs+3i3sT8K9GMqXZ1y5gRGiikBKAf7nrRkNQtWevhmBlbfu
nWHNnbp2BOUt1GNHTAGFutPlI5/yD+YSW4sPyGp6wXi/t91l92f3SrSrFU0FgJ61BfzkuZXy3sKA
snPkfsyxxTwEQGRUPnQbonSm5ASqWAjpBEY59rVIdlHcMzZg5BXVRFkrb/4XElueObArypvCtkQ7
9PqHQrCu9aHwo/KKHMtSn9qDSW6W06P81hlKYD2PKyjhix6APTs91k0jUlDZ2lWKKgZEz77TPqL2
4Zoa41Ad/JPh92YNoSAOE9FmzaZRj6MJI2zpAFJDw1FIyE6TSp23K+yfPthQY4l0ZPmKPEaKbDhV
0m6yuykgZEo+CFHLqoiUqRyD4hQpmtlPMz/0cjM4s6KSAsEtEqR3245wWQpMRea0wWNZuwdBvDFM
I26x8DzE/3n4PzACB8uHP5mJ0qfjMliaO/UF2uh+nksZrWwaMaa8HGB6rRbku3Y+CZ9+w04kw1Yb
gH8gtw82ByodwO1jkt2pytaqu8HBOAND/vYZ9rHk5CZ28RS97XxB7szV2TVPF4ARbuPkb+IkdtCp
NHa7dhIuf42Cty+dMdHpxdFjFKNilQGRQSNoVbhLQbDJ7y75P/iuzLhbB8k46+nwyfYzRPmr2NxY
uU/CTTgzjS391LzGc0U81vZrBlXWK5Pqx90e/g1YUdAfUlURBBPEcDfzBN/YhmV3AOtzxBQTd7/9
fvVH0Th1ObK1mHLDVJyJOGG0mDJ8Tk/Nk8bLM7Nd/DhEpYo1wmVcYn9+G4oIWHDbNUo3rqdjK5fj
oNmjquVbOshrAeJvv8HyVmVJ2Jx42Y4IzwOau3yKuHtBv2FEqK7U5NyOjhrfwZBxKCZM9I+V2nbX
L93lLzHt7ftCNcGqAQJqwRU7AGHLa5NMHC3xsSEfzRvTnfcrwq9SYbrqY0kvpTOTapytCAWuzsZO
MkFXx0bdfz+JyrkDqpyGQwABxfn/CS84p25TCB60fTogS6I0ri/nI9yF2gVRLsCHgXo7bmH++4IU
2awvWzRpQxUt1BExYEVUFzqoAjPBJMIIkuxL6VknVWKHqY8ZRa1TyVoJTwxQFLpCVxLNWA2sJPe3
YFpWc5JJJ7lKS8gHysQmeGkh2OyBuedWc+XD80dxiuvcK9FeQtyZE+cYEChnLCSjCbR7tdg5qBsU
ES2chRrTXfkAyHxt/gvCAHXkTw6xlErl5CbWbcKNFd0vMo3ydBKKKqM2tP14dclPYRQ823oPtbbm
3EMuHmnuHnjzCLINUDOprCX7+P+KnxNKKu54VSrrls85eMq2xoH0kUws2H6iOiOHc3JvaF6YA4iR
0hGB4BzTBvkBeJcof1ABVHDN3NJX1CIQQHn43fHWTGReQfOFInO4JZxb/IMr/L6PhBasCzvPyxqH
VjsFqFQpd8RRVx2ZWk+Q+S5XHiCpCIGvs3aCQ6Dzaogs0lh2bMX9uydEOCdNoPVXXi5Syy5IXVre
Q4y7sXd3C7hRsG19gbPoEGz3M+9Mt21Vk+nSX0XbnnvdAEBiYHaohLxikjb4jt7DkGaz2AcpRMyE
aoxvf2IfRlt3GXER+g2I55pojftGn+9eDmE6bECP2ZKqcgz1RcihPFrNDkRnqO4HB6O1W12ZWQ1r
CmLGQPzoy6sHUWlpcKkSsoXf+xzEnSV+h7FfdfIeiCM9c1POtVk4Sh0l+9uODh+Ymtmb9OW07S/A
EHKc2FEPokHgkAHRj+Cv6ZTL2P4/8C/9Z40yYCewi9NYp7f9+o8yF8WHYhhlYw5koWEThMYyy5Vx
ymKjuFkssBgPcmTvzxexR+TA2NyDBQIc8jrpkzpznBRQjbLuRh+BS9vzrJDhPR0KI/mlKKz4oWNC
LYn+z/OX3EXIM7WzmqWkCQ4qxMkrKx92Hldan9Nwz/Ugi6OLn7j6uWGmT52x+rVmVhT2sCyk/Kgj
gukaQSYXbegAnaq9XamR+9uOnCxRuNLwoh/X7lcHqijgcYnih2ndIKNgZfmOD8q9KqnslVbQTqPE
5wudN12D9FkiSkqBm77Ok1GaPQS0N9sQs/cwmtTXFsZLiSeEPItFojgAvYAJR6u04SCXUPZScooe
tXb3pmA6nzb83uCkE8/G0eoyo2143UTaxohkhua8Ofm+h4aXTkRQ+bzm3Z+8D1IxQtJogjXlHRaD
KKkwtJITKAhJvSjxPDoo1YO/goAfHPdKggubG7bZKiO+iSz9IoWEKWyRBkkZ4U5F8QmcK3kkZzfO
5I/unXv1pTiFE4XlJ8xlL6MJdq9+k3Cd/VS/sMkneVYtLaQNirz93JPblu+QnGe+/3ucvlf2TRi3
lyw0c6S+JA+HuWNcyIAxWY9fZhx2d2CgAaKVz88w/GFJx7yuqbM5qoXf45YAt9WtZGUHlDI2G6rk
/qEFIa/ywnyTxZWU6++ha8BjFz07UKhDS0TXvgxqXBkPsAygdJ24YcNtapcHy2T8bSUmqTSNfqfx
YCWBiax8NT2raDFkZp/TwW11dezO1AZxJGQIQDWwaDo806uZs518L2k9b2tfn5Df9SBQqX7cQbXj
kxNYgGLyCRy4+U2pDji/5tuFertHy5DDsBsAfuE6p7rS6pmVug86xeu7o1hhD6eVoqbwLG2Euxb4
E80mCDUP+XBiQWmcu9fV1nHW9ttdzu2A+z8f7qR4h7iVGymtJ8ZOIyciR6G/UWVQRNwuyneQCSRq
/KuKnU9+laT8DnBA930VcMh+VbgjgsQH+nRqSRuBRdoHubof718YRwV2JoYdvd/adT80PjVK7/Y5
5hI1MVMkWVQ+5Q/UtLT/I6Ua0G5YvtYWSoog1HsLBD/xtsuugIFg65Pr2UNBq9szIVlk+iWJLouT
Rizm131HovAGSqxli1vWrVLM+n0HY2Hlil5EoNPBVxYbqSFb/lIK8M/6oUPU24PxlClVS0+9K9QL
xomnOczek3C5fMUHG0SH7iKdjoHGoujngjwyhCYwqHDtRdafqDsBGPBBLB/Piqh1XCEfzCm+JqC0
X43x3ot5CQtI4U18nxAELX+dqaCNAhGXQ6EUlCB9IR/8CGzV/Nss7JqTgWGzdWU/sihQondnw38c
Eo9ulTrwYL9wTsXpGgVx3A0TONoc1gKT1qQPHXUeuRkTqLhH86HnMyWfrYjisy1BR4rnoViP9Pz1
oonZT53f1zPuL5x/e0K8MMROSsDVN9syEw4UJsGXe5tI+ZYDsTfiANYbO9oMiB2Iw1efrusYYi3p
v5plL7Dh81KKJ14v8j+WGyOnnSppMiPeN54Ch1MPTEb2TQRTxb2PknaActzTZCDxUlLU0RWk/2nW
7SJjf+lK5Qcl1NfOEPXcQnCJUB8iDqqbhXuMAlmq7fdzSQyU+lNIfLawBNMDjs7nHFV9odk0wf/5
pAx2/+NBWgWlTz27k/9gvLB91xG683aut5te3gVMTe3BfqDtydCr8FsKNmGg+9zDdBYEvKysv+bE
9BKwM7oAW/4n6d4hUlDC3hy1dGhSHGnPiCXJhvuc802m5wLEbKDv3aQ6PLrhpSUVOo3cutjYeXdE
movyHYhD56rgDWZULMYVHmXlM866Pg0QsdyyqrJ1yNLk9ktL17AH+SVluA69J07FczEucjB0UMF/
339RUQCu2/C8ZAFD0SuDRbQge+puh1otSUQlP5AB42+DRM1ikt2o/GFcSlRJXklfoFGphuT+o9OA
PwsAWhNNOIA7MSuLN+p1mP2g4QIZgLwJcsH+G5MjkdZbGuXpUU6JPEYgSZqazWBPSPY8nhuP3mZd
2Yxu1Zf05DaMBP83CM48kb1VZhCuYeKXybawpCSZiqW/2jWh8pKVe6Beml6W8Oey3uXrDdbu1byy
4VbFAW+dSUniWuSdGKNxvOBvEFkb2qb5r095fnymjRE+8oge7QTA7QCRfRuzZ85DXZ77SuarQ8aE
4Q8QoBd7QnY/GxvLOelXR+Gi88ovAtuMJD2nkrsY1c8aZSmfAHr4N6VPQS8cPDrc7w+o8ntfJrsR
PFTPT4JQbCVWxxH7q+Ba5ZTFu4exyIe9hB5sZ5Pr6v7BVQryT5hPxJMZZ3pgflLrY4VK92XqD2ap
iEqo2i5yDP7IxU36DO5huIMA04jglc+ohjD1dzyYNdkhTM6ZoLNArX3ZixYw4sSyNPabUMIpCOaB
o0EFE+BSsIAZ/X2lY04z3tlwiDf/4YUISTKIn/JfciwpqO+Br6vdy3Dvoxn0AisyvRfD5/IVLnVN
ysbTk+T4cBIfCxjlL2ezz3h3FbF1lvTFtHDAV/C3js3ykHg4FIjIcFUGb/BVlwxJhD1iAZH6YNp0
Tvrtm+e5Ap72u/tKmptmF3en5yC7dqKF5wvaHFfn7Dt9XYl0ObHu6UxlbJ4XxGBIaz4iT4naaWUA
4DOLNM7tff/FukYReXguiCZ8cNnab9gHQ7BVERX4S7THP/3jNpKH/IFRy1woYbrHAdk9+Hu2Ot7I
sfhbpDYF1M3+u/O46dc9+tsIvHEDW5ouEtsSwIPFAb+BMhXljQCqK30TR8eNqoyEfGlrTTMEhOry
eJN1imlbvGpMBQIIdwxawjFiZAbCsHM+mxwwoe3hgpcL7ZkCI79NgXOA5iucxmcy0A/MR3IjD0R3
70fpE7CH70MeZx9cHZdsxRGY43IemJVZMMh9qVosTF0mqU/jjuiC6VZuiJbQyPS4r0n3G049F1eM
VrfFyO6TLloK4vKcHmKY5eiwArGSqr+RphjCTtyxujoEDFy95esYvzF7xbDIKQP8bEVH9S1ffh3r
crrOcKbqR0/ElwSNHaBSiMS059XTNixxj9Xydtt0VR+0knAT8R90/9zxlhvZDwB1qQR6Ap+ujMJy
gm82eMnFhEZLC7gGsf/FPna6p1u/LYSZYqea7TWeVtFQ2e4IVJXjPrPCfy9/LBx86ILut8s7VWbq
zkuuZLoAdqWss67ZrE72R4eQagSnkOaJC/DbtYVdwWqKG4T4CVyoaGgbWiZmgtB7sxJbrTplDf9V
hr319nlj9pmmSddLdq875850Y8ENVWmfEHYKKXYYO0qJ0RlrUE/yqA6xle83c9MYyX16V9y442sR
yEsbft1VhtkEGLRiaoz8/4Lwtm8wsEgdVUPbnpu5A+EQhvKNWEd0BsnBjQ6WLk7fVYVTbpfmYH8e
766AdG5SxH1tV993D0pfgnIftMfcTaxFEcBSgBqLG0D7db58twCVIODDD9O3F1wUM1pzx+95Ypls
0sISHyIF8jV4Jift0S4M51TozpcIsYu0SZP4e4bdi/SBjZIexY8/zLcIkqiQufdXYT/avzKc+vvG
Jro3/GJYZ8VnccLFA2O8/Qpv49nXfiH/u9+mqhO8y6aJbvXp7hItdyuK9zqJst9FYCm3HqNBVFfr
yzcyFt+8xkLl6SZMV3Uo5xRiY3viM7Xm4KUh4x9dozI2zCYAfjGu2ZjI8UT2ILbhyVMICNBC0NSx
gNr4eepHI/r1WGBw8R30CMKLN+Z7uBK4zddesAWDrcZzYLQEMbshFqrqzUThATK9su+ggI2W7gGx
fE3OdXzEQTZY0RPEq/iOT1pn+7B+cynxZmx5v0DIft9lbPfzsqVNMaNYdOQh6frgcGrdPLaFcVRR
1W+SNfU7yWRv8Km5KDJBrb3Jb3XNWw+lzHipsYTaR7v8PWRoKdJVjhpEUt+/i6UfPLCyrOFbbnEn
XdUFXnMYABxb6p+oSCEIitrY/j79oTD57ScP5R/IPFA8OOVlFXrg7MkQnAzwdNSZYUPY58cE5P3l
hSJK81PmdAANpYeEJJP1acgPLQz6IvYTMQcLiNl0KSVifnvI6+wti4UwPcBWDHqkSfmxuwqa2ADg
iaC6bfIJPSqWnyT3qtamUd0w92elffnalOFXu4Udm2ml6RzuGfC2tut6jlJGCsk0/p7mymwAOZuN
2JummVgEiJeT6b88McqL6bg56MvHHgngC6Ua4hDAOwQRWTo4nFppuRy2gq0tIwT2cbY3VkaQk8TU
HNG6lPNvJapwsUl2JXJF6dhFEdO5VTORHEt8xoyUT0jP5bQ6F7T2tuPAstrBsb9hvl5SDWq+cfIj
UpOKvhl/ptM0t1UVly6iLdHfuycfrFFZu0RTwdJMLSsN9KEjkNyzqGHzCQ0SrWEiRpN3JKXx08DP
8qs5YablkdbuqZold+w0R0ummc1YdVX+/LqUhBv4e2pfSp0oHoClj4RxxhB+a8cNv7cCBWNcO4h1
1tAo9HUXaLR+FEWEHs56Q1iqFRV7WeHSA4dBJep+BuOwerofI4h59Qde1vY25obNmmhnmx9lY2Tg
kBm9RaTuNOl7ewN7An51cydDTDOslM1DR0BRQANYn5w3HkTKuXxQIj6H9kLegiHIeGzRTk5gfInZ
d150sHph9twS9gqgZXlFLVVS2KJ/383O10xAeTrhvrkZUyeTiPqVDmFzluW3VwZMt94HvD+iTm+Y
ngP4Wz3B1/5rHrOC83MjoXGNe3eVvahp4EzVW8rxcstJIuGYd6R2rXRVSw5KyWeKBMaT6GcaHkRW
fbSKnXf9p0T5waTjs3Mi4ZtA0G2c027Kgm4wWZaJVe+sbQyBx83MyvHBDJKGqmNzS63GxmQ+oZib
ZXttO4R5jyXoht0/DHoEgCURd/6opagghNWtCuF+JHbxL+Qw1RRDipzptlhBGR45qGrxg+ufvE5Y
T0yqeCzYWCb34FVZSdbGbBVeBd9nTKwyAIm+c6jmspRuYNALzl0XFBDfPhQ90zGoPXh+XFPkHEtH
Q9+8aBZCIhZPq23GPK46bNFVA9pNtzpEI+QXvXyNbb0KlGA2qRjpsn3XEKR7JuBM3Ty1p8ASWNnS
KxYpmfq0doCQOZ72fACTE1frdqr7k3Hmx6Ylvo0AR4p2A5mF+8tMrlygo+Xb6++scQxxFWuIZamB
H21cgv1NPQxD0BCDU7aQIGJCxj1rAXj6kAsHmtS5c57ywfBoCWQRlS98I+5/Yw8RTxu9/tCZfE0A
CSXCYewvlUsdKlCK1IJM84CllP7NvQS4B5Hxh1CF9A9tC4o0vRORrE3VxdAzRDya4cCG5hG1DavP
m4nDH0nky18hqSrAS5sLcB4ufKRmNiaUYMOWYHb6h7Xl5/CrwRtfaSEAbyc+wWbbVvEsMvYHp+dp
VdQ7NaKXbPsA9Oecw14HStFKdTZeOnTBOZ+Gri/VeW6qScyRiB9zaV1p3DzBvBpTF7cYZcacobqQ
4AMddTliS7Um/YR6uWGWowR6j9aU6matfUOaxydxYBMu73r8plSfXY4vI9g0Xm9koDhsNahS9PAY
csjMPVOEUnbvE6kaJRAJP+aNdp9+DZ5yrrLtevIbK5b/x3n0dEd/UKCKiGKJGJxQPKHa4fYQ0hbu
0/3XyxbjbEit0zbYNmsWlnMg3R2FedWBFAD/SXQdgvjgVzmiREHoKmNayz1yrlWqBKHdlSDQbnzP
TUAc50WnV6VORg6AU/Z0sm58E91+EpmYy27Z+lvm89FehWM5mlf/K4eNYM18/WEajG2MIHnjxCKE
GvyOkBYxVQDC0r+P4SRJzE7xYpXZfPCLKoSGPUJsLcJXtrMAGTRm0/NTv1NWAQj+7fWBFZiJaGxj
uD9Jwn0M+DPNwZJwPuu5266rnzCuVzBDXVSqC3EGZtbW542YeQzgnS/HGcVKc7fNSqa2jq6Wm3mI
Be6/gIGEzBo7HJy69Xe89NyzhEGTkjInG4KKqQIQz+q04lS8f82L3gAC69ssNpL7tmRtqfbjTpgi
wsnjwi0pvFsKwxqOH8DszIcBLuYzFj3niZo37m+YbobAtgkgY9S10si4K9DC4MCgo/9mnqpw6DJS
02xVYZcs4CCLq7YlDJsQpVn5AD6X/I2HVdlGrdBVpEWjeKIjFAP2dPX97X65tb1DLaJ/QCJqjF3U
c4iWKTMgkZaNJl4dRhT81xgEj+vjtMlNOMEZvKDLJGY/A1uNNkZ/nJBeCI1+Cuv+g1SeTKE++6uQ
RsQKqulD2/S7shsnIxhruMnRrZxzQtV8sCrsZMQKDNBoJ+RuHEvmEvlba91c33OEIPj7FnmYvK82
n66u/geKNi30frtjAi9LUXwCA7JJ1DoFPDyzLlSYcZCG5093WZmzPp3Fza4ZduZhH258zfqHJgny
rsHH6ASl+pwBvFjRD/Z8DshPLfMlIOFDckc2NSh/mHbrjINaMQYUqvWlKQt1Uoi9z/OSsnXlXzwB
lM64qMZZpSEXGRMUXEYN0Y/sjvljUY1JLX4c2L4BbaLu6R6VtosAuGTWANiuq6Lu/IQfesdH1R7j
VuX09MLc7yX3TDBVFJ0IZYbNi49xsgMoUJvTPpCrrt+GeGR5DXHx3db8QRduUBrQRzHDjfEMZrdj
972ja17n+T+OV0n3O/qgJPQ6a8/pkADfcHgI2BjacXQW/WKwkMD+EECmoqjbqQuEn9S6DVrA54h0
mJHGsTPIxEoRl2tuydgz1EJ/LUsvqm1ab6pmRXmOdMEgFznndfFwLvl7M8kzVLBbRE7/bYvO1GPy
t2+PwSTKhYdQz26rI0ky0/VfxJTpI6Gr/5qqiK+t51pKRZHhKE0aTdEiKp7UwwtdWphY4qra7r6F
zk1Cxr0rf9cD51UmDk4RfhRC4VO7HfEyr2udOHIC06Ts2YcpK0QPcqPw5HMcTRXwhYqQwPvdsNRE
1suSAuabmdBhH3T6DhwKu9Yi7sO0uYSfqdLl21W38L9DwtrB9Jb0gMVRriDL+b8IEAcbiO8b+w2y
OwuLuaPheaH7fHddjXEtnhlNJg3qW8Sbh+wqbQsqMxQmpz/otHDADW6bSVVPY6WV5gLzYFLnCm19
f0ysIGu2BtD2RpDWVaiez7oUvV+0Z0Xo83Nb1GiZM7Gu9wkICSq7XiosEWz/uIioe7DfkpwPeqRU
hISAJkEG30UPzgkdGrO/By3Zs1tkWzzbCawjh7CSSkKvypxe/jak16dScBANyb7q+roUpzJjHbBt
AQo63p/YUBNpsfxEvl9ig0zzaRhIQWF8QZy0ZTE+UFwaxY8CszieFG0mL7Ad4jZ1o7uwqRXj1rlN
Qgo8jrisIW2bW4fMWcqkVbo1oXakXmQL5l+Ao0IXvcYN79eABlTvNppVz1CH/b/R8XyUN237O57B
pLeSnK9QmiSZjlblUTLNGTqwv3tgvVjOfbBGwPX8Q78YOos30mBnSw2+r8eMLEMO9igh9sDae25M
Hoc3xZ1EsHGXu5Wkkg/UHGld02gUx/pkKvChU7Y+A94ytvRnRFiQESZ/iNenq3QcoDE4mZnkSPH6
m17AIASyhK2mbSjWrl+KXpG59LNDr3fMEmTNshhDpBp0XuqPMB1/Zhdfa5cqLfAybYxIfZSC4g0O
yPbV3rYA1JisCoL0TANuksHdAz++NM+5J/JGv1Ea93y68INefjIfReBb+QM7X14pTxR16NcEdvpG
9+S8rMBrJ2WQAioLDTeZKHQwP/zxygm3iA9rJdhV9fXmt/VvxM8eC4UwSF4GOijNtMhO3mKA26Dx
p9u2YvwY22gOJ/UKCm9G49Y9GJnQmLm6LxDsZUeaer8nbgCD47b+48OGRkjXiZ5s/HxFqqMImRIE
PwSgYHNUGCMZadU1/XFep3H03ZvikOgUkaEHt3p9bAkuc/sDthUzfkIhHU54QDa+S34xbrhgJ50a
ezx6f1zMofkAbhcdGxAY+RVXfeG2D/FcuJXjYKgQo8V7Rp/ECp5RK4e919Yxcnr7OQpyQ1tOJN12
PV1gs533vctxq8Gh/81hvNR11tDLLyQiBX5ep+wky2srxlvdLgnu50ZVznJT4wrtd9Z6lQhq9L9s
YFswaUI10jxV8FQbc++2lOEIqBHPXPuSIv1DtU2MWBGoKKKmRqB8du5gUKde44Ai1RhPG2towivK
1s0dSHakX9X1oaj9GT8YdUJOhV477avSw0E0OeZEhl5JbLBbtVstzuoRM69dtkvLuUzJJ/ypFfAw
nQK3TRMIdECl/4Bzq0O8r0a8a9xRl4XxKpKBkiTCPy30eoRrUA+LGrNnk/2qk/skh4fgQOUa9fIo
gZWgn7KGVqFkoNddFopzyrCGdrEABhZ5pZrJpz0rJuIPB7O/t5TaGSt5j3muChQrWYxkQ0kbxjW3
75XjwxQxgyPAqTJPNN+Aa076y/tCKmgyFMHwrPT0n3PpzPMh30HaFQMByYuAs54D6quZniKfvQzw
fk9nczQdymVkNYrPGmNch03oYkLOHpXa8X+zixDTuKrxGvKDVbSM+j0ZAUmjypox9pLEOhKNruQw
J6mycXJR9DWh76BEXg3+yaTNOnX9sLWIafWN8uegxdhB2NFHz32475DvppT9kEtNK63IUGxPF/DR
FkcxTnKSkfOyIpiPRWMKbQrs4X9ua5bC9OY/kHn/7AJlI4Zou3kZeXb/F8v08mFvouBtni/v0pFi
frzCwBDy8MKPfD3NfXAks5l6UUaudW+cX3mlducotUiVqGkr8GQ1Ikky3u1QNlSGwOy9sJW6CzcB
8Cgljq35sM/nY0/v9uDjaSRbntSL1kCTbrjJl0l4AU4loQdJkbclSfp0ccT/w2w6W1rTODrk+rBz
LAkivGhGx1Fl53GGuWLuqocax20lu/hnH0AQQnUs0o2tGPrNhPhbl6OOHaDteXvjofNk1bSkwDsG
30q+Au2cQXw/yenmCbCiTsWtDDcYXa04gPl4xCuUOJ9IxkP0vy18IdC33woi1DDsHyh068dMefGn
TJiAj5+Dc1BIMtNuBEx5SyAumL2slYMpR6Qvrf8jzbpcH+9iV4SOxAiZyvQGYRjmZLSJpABJzYsX
gD8Fd7x/l6iXAuM0Vd1EiHLquglWn7iAV8uZNcUjS3RfQWMEUBm7cOnxNqT5ZVXiFe8m8fLVOfBE
0ZE9ICMIdGaxzdG/96vL1qPy87om1sGFCNm+S+2MTSN0k1/Ur90d/M7XRZZ58GZAI86gSBPgPWy+
l8IC1xjmuPVqwOXv1z9dXAeVIWBLsNuMPOYkJjaBbQfiElvURoRDfuOUvyM3hKDQJ+3LIHXyyjQ9
d/EgJ8rVl2+QVdt1YkPiUgcZFGYu9Sjrfjf8YNrhMR0kkQy18gFTsgButoYM6T3JreTLsc8qsFfK
O97Rr5H6GVe+njrOwR5B4OMM0Dx9pnuzB5A3k8xz3Yxnvds4hvQT5cwHBx4lQsiIVlV/Ir56ePIu
u/ptyKTzt9rZxHsT5ZxJUoGylBFv2zWkxZFndpCvs2RJvk4/IDioRsTPA6yrHagnIUPmDJAzk7Vk
/Jx4z12cYeHX4S59CLwXdxpWQL7eoPf7bGRcsOIziE8FIk+FliJ+aaTU99W4fukLY5ylxRXeOW2X
093vJLDZFHicm6hbNsshM82FMeXjVRGNizUXzeeOKxLPoeJ00Gtd/5zWxkZhZrO6iIi1hGLxtK8W
wRGjoqCBo3PLZw1Xe0LVGbY09adwf65s5SpXz+cntO5uzJ/I6hTzbSe0SNTOxdFobq69WUcsJ/wJ
PBasy1gNdtcTdafaz8go2eRvIh131MP5O2BVOObL9YqWvvRjqZIwdVgWRQ/LpxgZMXxWIths9p2A
jdgV5kDxCCuWIhutmYFOtet82QyWIhkc3/IziBxwj7DPszaL5cGrV/bEl34pLgjx4BCcEOYDQYYT
bpkHN9tvMl/Q4j/JpZuQ8+HJ+b5lgEjTnN8vCgl6LLRUbtpqG2SBJFY1e/SB+ZJKS691ljSdrPk1
8AxGAHI0fBs+RLci29fg+IIqajN/cjQR/A7reqbKJJTvpyayOJ6cgfUMEt4SJXQkM4t6qDaIi1bG
+VLEakeHl62QDo2sAutLyjldCzFp1iGX6KZEZeMI2SyFnC5h7UDofSwq2xLJ7cfymH/7/7oF75ya
6xuHlcd1WPTZ0qSaerwi9R1H1/Ii4c82mcRnc3/VUdW55hHoUnPyOIuHTD6Mfpjsw6ZO8C/bmjhE
BufmS1qe7L9HkTZS+0fHPcmO6EDP1y/QH3mQOeBKs18D3h19FiNaEz4SVsov0fxGseqTgAdMTmRH
AB6TSInoM0AfQEAThRApoZLh22Fb3247vNN4Sqt280q43DaIN6wPhAOFG3pFv9m0YsdDD91qC4q9
T4JdyiWBM/7vjfVhNf8cBfuJZ3QM15rZTslvN0Zesz+dnrxLWnNbqcVsMJeD3EOxA/LyW/DcZNKx
61uz2WJfXXvp6ocyX8wrvr5+CU8K0KcOflD0dw1wUICy+6xiPVun9m0MvM1v1po6/bvK4sFDvg1W
+jU1awxN/vgFSJj1vlDNIiWcXl6JT5d0NsxnJl3jtIsFI7X7oHeM+40Fu0jd3xxjb7Hn2XtQAznq
cmRGi2cKUrtonyMthXTj/UYWRAv5lHLsc5hx7RgSNEXJzmw/3/ce0DCvh3VDqMuHn/rWVyPVYLHY
fUoG5tsmk1PUIa+KUOzlKtnQYAT9PaD4aiNgTc2u6HHuq2BrQSj9NxzfwKEUMXJHP6okK52LhCNV
hADoPzAREoibgJ+WjrOBjr0kqbpUF1Eks2QZ42IaPjn8MyvDTt0edqxNl0f/tL8G/DsdRcM+GzVs
+tk+GGhMuBVDyhEjTviJRhGu6Jotf9oGrXgyv1lnW/kfWWhJKsTWK47Lkbwgaz3Nr0Mx1vYdLBnx
14OfEhrTEFrRKu8xlQAn6kZQ1w2nZmO4P8tVFjt1dtZjG8+wqCBQiv/gm4kc+90I3QcxKpUFbkSp
rJHIztAoT7+1FbzRry7nsnBOhbzuwmFT6QcWsbsSkNsxdYKob/qnknNDxdEA6ClGn42yC/OdBJg1
JWjvhqccECuZQsTz0x2QlHd77aPXjTRcGyML/mM0659q+jViX9woCOI8JNtJZF+a5Z34C70Gch52
UWOHHQu7/8h2S3nXvE8ReVb52HfGK+wE6sP83znciFZTPTWOWK3pl+TYgKLzAEZWrqDmdD7dUPQ1
TsUdUI7/B2QRFino7sMWGx/doKdF/AGybdLhHMwAw6Yj7dBHuUCj8pbrtjkVSyXO5PyQ+LhkEbKA
DOjAoZ23yO3YleUZDtIAkhuEDa3T89QaRyhD05BIycV0kT43ZgM03r9BrYi7XLkCdeqFJ3eyK63x
8f047INcKGCvLnt1rcGSgoOgut0HYZYeCGJ9tAbnBLdeXbD5VsxrMcKxfEQaBd7sJCQRRKURqS6F
oJpAV7dfcwVsjIuIDNYteEmdwT9t/f+Rjzgn+JHiTG64ZqJzbPE2OSTCo7jxCqr1W+gXPovdR/bz
Voz6TosKYFxWoqap5tKLvleVPp+QEd6xV3xO5Tx0Vt4bCYZowJdfQ82i0UiDhZQNzzgcVIgowYq2
3z0wlyvidP42/4lCqw1XOOsCtNfhWVWwzbjYDbt49OaNwVUdyKsPW6br56z20N8qPUo3yQxpeW19
9rmmOlNfWKyHwZqtfj6V1jd8g4h8oFKgEWxh8hy+8LvpNSl6P4WvJRoDdZBZNIQDPrEyqfojBvij
NvcvaCm/bV1g925GSdNCP7hRlZNta1kAr5zFPAMXzbl23xeZSY3MYPTYXUL1M5IGftSgSOnbOEWg
Zw0iBFL+BXrPSmcYyP7U4LLdI/W05iHKHPDtuVGk52ZI4NOfiL233/7n84LRof88fIL/MTy+d2Y0
JgUhmBmn1xoA8r0H5Gc1ezZlDc3y7ieBqi6F4di0xryAae8sB8LuFmZfNGxb+vYzJgr/FbBQA7eu
mOWRIgIH8JbTPDxoRJHdVypW3oatCq5gu6NiCn51ksUmxcTMS7KjkMfvlMMb6jSt2g4oa73C+gbn
iglF4jqxYV6Synzjt38wxOQsqlbxKdnFGAEHOPc3ub9+eoHG5GN+cYvhx40JSxwytC/OxsRUSdhW
2257xs4vqN12YitWP/VMTae7qeg04hNcxw2yWCs/Io8jZaVbwFTKT7/2xHV2/TxpqXrwSiL+lQj5
TXPzZb31TPzkUmv/owQ/585udcwGqOrOMd4jiX7FFTKZlieuEtPUNm9BlHGChf6HwgoqmNYyjPyW
qelw4QItyhhu4D2GgCD/QUCUPRvixcQKzA7iLIbdPe5p6X9bU0c7MVAXT15a7NDBOLTzQhrx5Ckv
USzcnBb2CpPm89pGWU7keCDFtkKgU1MIb9yGuyLmRTILKtusmp+kM4SkvKK49ZTQsfroh4nmPVUg
JLI9Gam8lfAojwy1tsxoYvJVoLpAWqmcLx2LfzZywnfXmKzwZY7GMeb2Qov/JFNQuPvO37Lu+TYV
RZKMkt3VfBANf9ZSMBK/czyJVggLPXo+EylMv5KLNVxeQDZPaQ6282q0crHKbyE2Ldt49RVp23I4
UioUGjezfvjnReSl6SF44mem4ykihK+J0IRQ2tm39QPneee6fFG4XHuQ3e3W7l1HrexAk4apEEK1
1WIm4doH1BilvlSnFVwE4QgfWsAZquzAMBwkGBnaURv8n4+kb2Q98dR8fSQ8+8lONwF7uhH1ABNN
6R2SIHzTkD5o4WOISFIsODo+D/bTnR97UvLUzITZOY9sQj/49D5TwuxVz4YWe/QRzBEg2YiN6N5B
jvD4nJ8KQpc5I/HrO+fVQzUZaBb40XgwVFmaDj601WztF0qUwlWJM4lKFJJORvDqYDrrY7QtI8to
wcEWy6aYmfKWG5ie0/GzhTsb5GRq61OSCxJ1xhmudvMn5vcA6GNYYxHU+Tv5bcbn1HjYkIqsCFqq
J1gMoNfwiOEepXdwL5qRrmFQLgsJySzXyfmC44EOhCx2LvLYF/KbWQ4qc1H6FZI8wgOt+XLNLl4g
ylhfjAnE4ic5b8eXJKe1OPVCZxiljVNIH4VCSKobdvUpbzBWd25ExugP6dO3JkCmhiQ6lqTml148
0FMtyogasMbzwx+HYvGAYbJwJj9bh1EyoUdKo7KrKeeH1sqY3clYMTq/aw62/PgnbsLXYItS1S9D
mVQEE8fIdCi5SzJUo0NpdDBvEf8Akz+/BqhBCyNVMl5x9xtaPnhiEny/UOZfIb4JCUCsJ3qgCVPY
xEjd7CdhWaDPYg+i6bivjUxBFwoexVrbElGgwOSiH7c8Fwn0i8lPwH9Mh2RGGEsdrCk2x0Lgc7FU
5EkL6reDZhJ4wSdVu5GXpEmM9RUYrv9iLpCGp4Btb0oVOxY4yLhccEu+EmdQzMR9rJhkzpt+8aPQ
EWsv/thrWYWjj0pLq9E5037H4z/CVugeDHCmtXcVx39mZ6NetjWcSqEFUS321ud2bve1/nrHNLSl
tmAiIA3u5MRAlDUisWg3anAkQhcxksRSTWaY+mD8Qj7VgO3SKwdwe2TnNZiEsW3ij5gF3WfeRm2l
kB1TglzmyadQhXinLj5JiPBd81HaGCy2mBSn3rNunUIJ6ntLwdXkICnYxuwJQYO7CXDqkpGB0U2e
53mT2vckzvcS1AyxWoiWtsmMITwcdrv/YP+PE4cU2RGrs0xbafTY7b1SrhjrZJO1UEjmeFgQTj1Q
4vrrhji/lutVCYd8qkuVyMenGVhqyMtY4P5UqqfpkJ4Na1kaP+ENNrWMTyULyowu0FyvTD/95mLr
7kDVgAKYXr3lsG4ZHa+mEHL4h3JBCT2rlyYjxHJu+qz0h1T6UqEqOiTm6ye+VfJoEfxgqlNIfqI2
rBGZ0QW4KgU0NZGu2nDXHqi1rHiid0aoOB/iMT8ecdQgml4BPRjh+ksXbHpKf3RlsD9TYVWESM3+
ZKDsXfR61cS87WboDsDAYItCRMC/WE9uIFzo7IZBNOUU2L/VBco2jFp4ZZr+qot/J+U8yrydZ7c+
ohCYwFteMZ3TRT/G8KTmDoqFybMzbDvgy+Tu5xLy9L9al/QUGjs7LciCKKp8HIW2Sk+mi04vdAvo
2OJN3HOMhTjBhaO1hrNTY3bSMB0uf0RJbahKTopnQNW1pLWz75rhMr98R5R6Oqy3ioNuNqrWAZCs
7XJTdeNv0kPkMuReqn0SY3e88f5YAp96hG1LKfAzwqsnWPBefS28cutx6sxW+FzUNSvkQGYFMt7B
U4kRrrq9iEDHZ/ZYKnl5GryY5Mg2KTKP6588E4s/nabavsEKpEervU4aHCJKe0ZcLiIyExJpSXXu
y1/4wXQ6YQC2hDpoPYGqAuZKstNyMptjaIPk665hFOxByuOaT5Xl4xbSvgqO3SJggpR35XKLnWSM
SP5p4NXUmVousWM7FEjA1PtoLH0+kk6cZFnybzy95ILXgY2D5YMjVnpaTIekrGU7ePVhQHgJlDdp
X58j+qep9MjcSwORwYW+ZtbpADj0capYJNcsqOGaZEugkMa5wAsGVrEhn4wwxVMRB3bhp+EZQndY
lNZNd3hFcVgOyhxLjXwRJkLPk3cdQG9ONgcF8orgDrE0z2TcV8kzzabFUexINVPZY4Dm1bcgohzP
K7utnqqsjB/mX/V1jIi1/W1N/yVwCYNoXpR5bM6axY6BYFp3sb/ZN112r6sjcTJ6j1sbJhPIUXNS
RFUJJQi7U5JDNnH+BpGocibb7T3zglyfqkqlq4gUwAyyDCs9jgG7vWeS62Tou/JhBOBp5mJ9vVsu
ZbcjQvul7Ea620t7sD95G35UwElSg2r+E49FqrVGqGmij16WdSAv4zm0cA+xtrZ0Jn3xrCFZDiCi
1gO5dVDnH3axgz6ITEZe83cDIwfr/I0nJuzAPF+qO1NweVWY3oiJDEjj/CMhR8F81XMa4w3OJBIP
7ORhPZuDCK/4q5b/leGfxBWBhvUWnuWbCTg0swhzEeMJyxomrAk7Iq5bKckg0CrMmjlJpNkLo8r9
TR07xV6UQ818n0caoELkbLmcnrkf98CESSYuiGPZ+ogCBmW+btjlF+GBytBnKg5ZdBoZxFBmzrP6
fGAB04Mj7jse81pay8vWvEgO4mF+U2VVPh6UarmNdXrbnVL7iXzpuIfl1szSiYlacoA81yWuDMUt
+hldTsBnlsfkqtrbJh7KT/re7upl97QwWxj57Cr/AqSJFp34nbYCpVXTVcxVE4+uCKcKnQgdl8lF
BDRM/lNrQB9zPM6j2cY9YIMtAjM9z0og4nYv75QRlNWMUg0qGPiM68OtU8vfe+KMHd/OwZ1K8sXJ
livkXhq0s1PDs7zaWUTNRG843KGhPz1Yy6xRN2q+XOJOLybXgV/xvP3wQZYHRxVKPGXVvft+XVID
rsiFpid+LHBy1KP2e+CtlX1Ar1DXyMwda4sriPcuU1RNMz0c53eD3JNj1PMvbpvIql3k0FJ4hFxU
av5XDaFYO4vDNUxi6Tr0mDVe6jDNQCx9GoKXHq3A/GtS45hp4LAbP0wnoEVYIy09d+q2+Cnj8yto
ohRuZfj5l6VgFkEJmNorQycO5sa5I+eRpuKdeGMRvou9FexFaXCovSRuJYHq7ebBaQ+D2Yz5YXIs
RLmTaRcc38Anaqkj6SZRcq9HLHgx2bAuR8TAy6/0CBRli7NidcN0CZ/2/bKHCAO7rDQ0z+Xz14hp
g30cAfEJLOEQmBp+kAJKGlJdsfe7dfrXbCYxSIcY47ftx0M7F/U2F5GgZwfSEPKkeAu/v+h9RhJ7
JOw2xTruniyBPtoxRBP/x20pf0FaxqHWIjEfQBUEwiZaUjdV5ME8dO4u2m9Rs6BeysXHD5k8sVRI
8or4a007Aw/PhSzgPBtTcFAHXoPIKHOryB/0WOU07DtEOE/0mzYfenrd5Bpc1XIhn6FZ/F9l6gd9
r/JcHPh8M2tQ6p9iWLJrtikmxAuRxrTdjGK3T9JByc1cjEdnJyLAaIe36YoR3qyHQDsvPXEyKPqQ
81TBg/zzCO8TlQiAvYGNlHmjSewgnDCyJ68D+feleJRvtLiv1QTo3ZaQTSZOe1jnwVJeMg4Dgl7z
tm2glpXlWwcC4GDlMbtFnY9RJzXTjOUCj8HpBnAm8+cX3cjjQ+9LnPyXTAC5KIUL/P91CyCoqegt
VEhYejCBaBwXcLgwF+fSmH47KXvE+DEz7tGWgwfKLyte4YSDDlDbtf05iQG0pQV3B9fYWZA6C0Z2
RL+P8jCF/Jgz/J2ZCMTIKS6piW9syT48lrPWxB/aslTJVJf5L0leBUZNsHvJu1EH0i7vGAk68bZA
foIB+k5MV9905kcnTgqTz/bQrVjxScLA4rdNfIT6f2XmfSYVmntJYmfitjiL/TaQZBDotImEzEmi
3hz5x/yfKIWuURiGvCYKWIpxSNqJGnvoIQn1Nk8hErZc5YkQ6zb39ujwKAVigmNETAfibFq8YmqA
MEPYv0b/F2lTloCF9kgUlXAY4XUpJI13EmgIk6+ureR3nOGHzG/h00oguKtQhseKpS/qovP6Uoqm
CK4mSPByz2oOa+5Ns77RjMBqtA9R2C/ZWUFV/O3MUzMmaUEoP5+dgqSdRYllNEGBx9X+lWS+BquT
ejJ+jGl3lYrTHnUq1VBWdNSJTmci0KIlYbDJ4Yr7x/UcYMo7kDjEZpnCIElzDn50RnMjFTwDGOg3
iykMyaqknUST9exSXO8d1f9JfjQ4IJ8NhMaZiEScdpUX+ym+ouj2wjv0Ha0qYZh/a5UAHGg14fnP
rUEbX+JtocNgS3hXhY/UbiapT/9RX5vDIGYtBMgp//REzTjk7DRqasD+ewleLwoD41rvBO2QV+Zj
5jMQN67iIXHgXnu7kek3FBrsSkkZDQOm64KGenlAdtHHeXYpVCHGM5xaKhilDZed2qvLSpTct5Kd
+em8GfSwisqtS6FfV8OADD1RQfPXCS1XLpxIolFP7f7odyW55kEQe1JxyENGhgbuVdxcgEQ3oCp0
aHwf132YQR7/z+7NdTqLR1npGv4Z5pJAMG/ixOCSNdRqw9l+26+G2Tgmao9Lyq8Xt4FRDsjMjtad
PIhJBe6TWOdhSAmO9xGoAPEHUmONkxOfWt9/e/QP3GQkUPvl6DX4OYdqZzCq8QNa0brBHNpNGnCS
AE0u7oj2OJCa/NgJfdTa9HbWDhHqUAHBrNw/PGFzbE9siRuJSIcmOBOp4LnuzLNghERoO/CMtIcB
H41Qs9Y0ljY/wzr6uE/L5MMqFYvzBjS6K3HXDs/zHlxsji8NYIN6zC39e/x/nYQb1efIGrLjYOyZ
h4+dm6a1PJ6rex0Oioh06Xpz7k753cT/H5wsW34OYsAfS2IQ+KvFMI62D6MI+CiRusF3Fi8UikF9
7bLLhiqY1fbXtIj6otlq0Zqr2EQV7U51mxC2jeiK3AixiJUXcc6G165PppAiCyYpwnlp0kC27Ehi
J/f3Hx9P/UqSqS3xbK6OVGuLM1UJBFbmePQ773gXyPP/ImTLEWp1rLL4oo7fGloWy8XzM2wFsazs
6K5TW0Vq9K81gAfE9y09JCT6rCioG3whqG/ZoHda3dn0KKpeiO/Kk3NgaHe8skKFWS3F+sBlsF2+
JWXntOYqW5Kcs8veQIu5HoEsrc46n1R9gqA4glm+Lm5yBHniyaIw1OkrfBWxTbVJgRtq9kc6iPkT
pOGyxs32lCBWOqwKalNF6rB4D00TBiy34CWj2I9Cq9iNCg6B11eIIlSHEjtCNpFeE13c3fUkTu2m
XjgfcKu7LHe+W93RGxCs7bCtDXkaETNqmXjlb+mkufFqm56Fd1EBrbFpamgFEYgH17cIgZWLdmg5
3fJBgsdqoAHbrT7o27gVjp+p55gUH8QgUBpXT77QT0t4L3m9/EIKatVpxPiEKN73r4T+TltVEcw5
/0T42XKDkMR+etsGfq1ijCPoijnfTddqpr9de9xL7hzMkSTV1Gc5h69wyfIphYXC1crVM84rGyaa
+WX4Z8sxrjgupcz3zGGWeWU3dVHJaYRCkj7wey1hkA0KiAUZe0NS+rb82UVaSqBqC/y/URx1wOnj
zuT7+amGSHm6TyBH7Ewd6uEObK5DwQDiwOfDV0lhlegw1d3GqK833ui2vCxWkfDYAju32G9Il4C3
yWaUVQWWZxALp/z4Uj1ayt96XKxoIr4obevsD+Xt2zsl+X48mdR4SA2IrketUDryzKChZFjxWN6T
GZ1oCbKx0m0uCSUK2QoQv2lUPsM3wS18VDKnR7XH1zbnDRUVnb3KDz1naAaO/CYlfpUxJ+FjH7Gp
VIkL0pChYSk4dQp9iUkNlVRiiUll1aZNzorjvC/LH6ikXjoE+QolR6kFJAA3b1Bd4FlCpcCZAlum
/M9etUopiuIst9Ku9y0ScqPWn8a2UszYFPJ3bMU1h3K4KG6BOXd1P69P72gmgsymJr91O0IlqAfY
eIyhophjqmbsKUKs06Ln/g32HIeZ78DSxIXSEP8ODQhg40lEzWrbvzFP/+ReI5pUypc8b07EK+5D
iBSM8nfW8sHrOU2pWS/hELCBQgEbQckUC4rFi36aWNRSHIYjl2958+5JwdDOyiDKEQTDRxAmCvKE
Qois/7STb4vyiMvkn3TY419V8jDzV97ivFuhDFVDxz20whWarXpMFtOfonVnCj7X586Dx0PRtwKW
59yNfnUNzAH8zvpL096gnt6woN7Qm+xCyUmSm2k0cGBV+PRh8Hyl8ebv9Qikdxlni+En3LPVu+lN
6Ysgdl7rzVB+IN7zXSYb/sZ1Gyt5h2qhLZOW8hT8cVG48IcfjGYX0l+THthKCZvK4iL1bLjl+jwG
Jd3ceDnmKJVVWvOSbbzdGA6gxgsIdCNHh/SLia2tsba21oQxh9e5C4YOiG+lb/MNpdXNnxONVelt
5bmos86bSdMc+9pPJ1JF7TVypGir8MBiSVRcnHctE8B59rDyPkREdtVXE4klevmicSVbrQzxYLyO
lMaTEJYuh2Sj1pV5gtCCc7YZgVo5LC6ywCNrYMYSj9NJj6+4FlXMfCBGTtXg4Gnx8cyE4a5YuaFU
zxuvthwkPaOrvF2/tPdffeerOVrhmFsxh7idQJkt5TfsUEYyZzCrF+rGxr7F4lnl5RYzWP7eylHa
Ze8kUDxW8AhXiNlLVoSVqKO8AD4A+my2HiF/NgXRLIeVWCC7QS85q9TH6BdCBYg328utbgrUqRcO
CVSWu9R/SnNgGZAUifhTTrZ8mULZ8daTxJ5CPu5Ui3mZW3Yo2fHwraS+nfTVcOQTAPHuXKoN31Vg
SXhcyEW+V7JLhGS1q/DaeVFJGHv1yCp0VNfvZkS9oLCuobFnh5OSRY8PMc8BJSC6DNkE/LRzMNq0
Tayj91hOb+U6GJPnvZOXv066X5l6Ev6i8iwBaLREsTJkaitoEf+1GCYNicyoHC9vdKKUz4VYjJN2
VuxZob0MRtJBm27KpMB/ABBO03r3C+xQMk3/J6ZwCRf4uyajytb+lrEcfnHIMjd8DbKcMGNbwWC9
3yk6yXe0o8SWc3JvdZbyLoYtZsk5wqwsCe979gT/2OwqV7onfQO+QXuoZhdkIUPXCnNgd0HYRP0k
ebPhsHJZLkUv5/5jQwCwFwJfFp32jHCuVrPsl7Pbzqnfkjxws5PtgACJZdrkEuB/VC2iqVZEwZwS
zpWFX23Och9Y9FKRg5qJ3H54AQ6fUna5KNUJcYix0EiRW0T//+aTetD9Vrlb4cgJxJ6Y0PfvuL+W
h0A5xn6VsxUfc6K5iX9c3k0Omy8ruuSyEqCEaYgB/jIsnfeJpLcasofDu5hbpc47BPYEzwGo7+cd
58BFxMpXa5c0vTMePCj2mC572K3mTwVDqKTJycv5txSbfYeyrLfAAbYVEw4hzSrRbGv5ruycaHKr
bLjCLq6bkS56Xl5EdH0D7OZlFyPGi9dots7f1QdAEFjIL6fXFtMkP22LNR0J4XuNYJE00rJ7jfWq
aBHYJflMrPRl86+tpTcU4YQM24dHRpYnIi/hnetUdWkkO0s37QbOo0c52GdwY4P4f5sKvMUPKWGp
qG+CK0GB1PDl/oKxTaetvOtB/Zi9Se2iHu5VJDvDkBsKdeK7fDTqeTBPCjayS1pxauoFhIKNXNHN
WmpGAvOVlq980kUmT8DOg3+1Lt91Plzv9V1f3IjUTowo7l+eGDfgMKH/KTL+INRk9KaoseTS6tkJ
fEygPhysnB+ot2gUXDAs1yvf2YwHrtTQ4u64rTQNkDoFqvpOTGEdXf3nZFlxiQtTRP0P1KCXuR+I
wllcWKjUDDqVHOGTgGBVVuRM1vk6wklP6Kc7ai1SXw+5JVJi6fS9OtK4DlqZZ3RqIMpCuk1PnGFy
qpT3FSmTGQwNeHLRGsSAjTbqvQj5kp5qkXzYOjarjt2O/2NA5Eu38u2bZZscGbBmhgvVY0aJED6n
mbihwcWuaLq0YgevfMnpenYtY2pl2HuccP538+PsXBr6Cn/RX/FsAVrZebrRFT4JrRklrt9Eeuwc
aRtecffykICyJEMNbYutzrOrpCKV4yqVya9i+//o1Yis8NZjP0+r3pndASKtm2EE3I8Ss2yoqY3O
vbsOxNyRkbqBYQVEYIccbMDXdPQ3HWXB3y3RLObxtPmbSwb11vMBiPiYZgbftzUByZHBf9J1qe+U
4oBesvgUNeEK5bUTLoZwc3hK5PN1BqmAYh9KKZBsJByaweBvejw1ikbEZAHaNa4Lq4RMdF5weCue
hHhPKzKaWefbc7HfVCFsfu+UQkux6OY5DDqY+SjA6AcQiKRPVWCPGw8kd99fZtVpCZ+OS0NLr89v
MkI5vd3lkwow9YBLFm3Mk2UwshIL40xl1t/6wwfyErBfSQUYJYw4lZMu3u/YG1G8uy2HwLYJMTA+
XmIP4gBegysaAldCQk6r02dUx/2NWfNrjnD6J5auRWb2ly382wIScdjKQp4Sm2tm+UVa8CIPND3k
R5k1kdOLqWZxJ6GNDVdFEw1lQvaYnHr66pYkzFLiCkUUpQ2y4L+SK674FT9q2GwoQ/pfu1kFh7ni
eq/PFHL4A9+823reOYJ7bHsJTTYvrsnkdS1FvfNO6C1UcwiDgjXYdo9eCTf1wBgYpGXUdApNUggg
dLdGmhR/I9WWqBiF95YL0E89i1Y8JYFcAPt/1N2wcKFgTbdLXCCJD9mrw6VfsKeyIuvzj/tBOxW7
TtAM/ln27nmpJgfIakmmoZknNlR429Gq8akeBkyI2gyM4j003iamS4FVH85QQvPLBNqyW4xCGzL3
caVkr81bOfXB525R3KwjBRMmKuDicy+GRgFfJEVut03jkMezw6Luu5KcwsYNvNjYk5ch5hZJXusj
xgxiuTkkDT4OuV3bvyLORFqntZ0oq4UXnTbe1nQ6D1WcxruEpppE0irrIGwL5zgrBW4bOxtaDPBc
7Bc04Ha/PvUAUh9fgZkHFnv5f28wiXci9Uvge9ZJkjXjY9zixRm9HgoFpILb9/PeWFHR8QnJyhoi
owQph+q9mkVZ/wh+MEcpQuL0lJsWGgEWHCJTT+gIQ4pY5myqbM8Hv1siMcJYfNCbc1g7H4DACfBH
D7O4gGw6ZkWVRXZEvggLJppUz1a91zPvqKPf8jKB1XOwtZXLt56P3SHGOowA4V6lex4WyhuI/uMz
Dl5NWd+bL2j/aGQid6G7c+1sdOgE5tvgMzy634nKXo3FXeoYk3Cf709wcQcMopQvL9b3Xeh3HQg5
BdSWI1Al3TSj2bmxAVdaLoemb9x2kryl7ln38idYYF4p7zNwsvAo8m6qpv+r7a7fPD2sv8Iqd9K3
wL3LHKtHcKpbpfareSGPIWAuSgYZDW4a2+Lk7jf1J78VveSmLzFQu4M/NnXo5zVtOoxvEIkF8OXf
0SxUVWQKoXmYD1seWBY+WcCxKSyKsENvOupOAs59Wa22OcsSRP1XJqPeGs9Yu3vHQSp0iauQICq0
YgT20ZYvoapJc05f2S5gZJAUzBK12QGf2GIrJpCI2jigBwgtaVfYxOI27YwuQWgZdBg0z1+foNge
1nrn2n9mf9x5Kcrgd3u6AiDbANtmJ9wGKv9yhuCJs566MT6QJjnJj9d69L2vcWqQcFI391PTl7vG
wnh2lJ1iOj0M9aYmsUtHzkKsHs4oypQ+9zuwOtPn3ZBd7t+LasiSueBvu2iiZIR3eTreSDZ/FcnE
bHWlODLyX/ZTMopsejVB/UuahwtOhrkB+p1VcLksyqIEqZBoYLHIbVeLoptUtKU2LcpcDCJJ0rmf
pzytx0CZVkhExdVydziIMoUsG+TtWzBKYBPUat+lk090xsD7ra/+dejBMGRI/gbHxtotQrKWrhf7
17pyyFRJsAhLdEWad/awN4yN/xZKGnsDgM5NUA+ctq0ernzELNoUi/ZDX1l7zqPzUDcySyjxKYhX
RnUYiNkMvlZ49Kslzr5Sm+QgaxZgosIWbv16A0W56TA4UM5+1XmD+u4cvyURDtYXcVA5dRjtNgMo
k+mPylvKqEbyjKGl+Dr+p+YHYbPRexIUXhICMbB1ndyOrBJI1I60Zew6iRa3TWU2RaSohYGh0dJD
MoabHTVlOjO8F2YcMRaAFL+SA7ymp+NWcR2EPm68iAhNm14cR4wngjUiD9wPskQ9O49RJIzxqT5b
CY7G+KwmmNJTBhPYzbnO+GGpVLsrUIDljFw/XQ5f3+THUCJZP4HE1MbDqKIo2MQzjaoSj6ls9HWs
gA2niByD2edtGCyRbUa7awR5kFW84Mt3BA1ZGSmRBCO0i5BmiR8iAfodo9Ubzu8n/ZQLJ15sjk6s
VCAjhdLuo2KRjsTShqJ3Z3su+hIoJJufR66r4juf2bmCn7KWaglBTIjiOmH1V7Pa3AhIqj9WxaXy
6YL15u895tCYG7vgAtgONjB9vOFGDseAOMrMqShu6uiXUU1GuYutHZ48EQmoZOE3xC/926ItCRYH
cqt1fLD7YEeAqzAutyKYHYhLNYzpb/yWV8qJ4n/rWb5/XklrKJ60G8YFVeUIVBsxYfJzC71mO4Lm
vUrXDKC1y9yt8NY5v9aXfrC9q+6WuhHMFkNQbY1yEnaqw81IuAqJyF7DxVe0c8pp+MQDiyu9nQ/+
0KzhCD5RYBlpl+4NnVkHnwopubgatvE0Pj54z7fNJJdB/HDJlg50wgnxg1Zrb6PyEX+gRwYv/fS1
M32vKwJDzoThi/1+G9O5Jkekujg9C30ZyVzGKv6h3YCFJYS8uQHVYhgFG62gaIlC3pa4tBP4H3Uq
1EUOG9xebF0PDy0uv1BNuoXp26PV8YJry65ImUVc6Y3dhSEs9smF5Oq9uAEyw6Xm7MuEVNOltF2G
q58shcoHoh/4g5TlqCp+tJvPLCBDJG0QD7PrTQc8oM+KlvM7RVAhOLhRkFXEw7ppjaIXHz1WDin3
4DCl6DqAPHa8SMkqeQ4ixZK04hukhwj7rgYIocrV/5LfIfjszR4H7pyM9W2EHFQnNrFGdXna7J46
0fBXVUADv4uJ24+6DCnXB75MyJW6Xo5B/u7p6XlNQCY5fjyc5EXTeKrXH9nLrFS88X4X5PxclIrw
rulD0trNHwgtGDcjKhKt2o5RQf/1uQarsP8R32baejuwhwtZuLsrZgpFng7hLwBMiFU5Q5neHVqg
J31SuvmZteEdzyXeGpymjIWeuvmyde+npvzKQMbf7LmfD0t/R4fabHLCN0yTP8x7RRAgAWSn5B1v
S6uBxvpuUpJzAbjIMoMiC6n+2XhGdu6rtwy9fnB2UYuhsc1AJsCOJjkyH5Bhi32CYM9FoeZWaotd
lQHTX1QJ1LcE8Xzdl/ag+UkcSu34OKgQqy2ExpXdxmIplocwo8Svl8WtQqjB1r1MD9oTOuZMO6Cs
B49Zo4S0H4CQPQLSGqOXgtxHIPn+zte4XdgLZRS6s+A/KB+u+uMsa/4WMLj5AVAyVIRskQTxqXJ7
eJo+Gxiw5oXy8/7J1SVLcUnT3A7qFUQB0nP9vFJi0kUA31HIkQ/KS8DTbf3phXaQsMmh/UnqKCm+
ok/dJArStJs2cIexPGpdOGOWJfVAYA1ANIm0I7y6Nt4EYqgQAmbcm7fo1UZF7Gqe0tEzWeh9hS4L
XlBZMC0B25aCiiHWaZUNuhprpD+hCGIWc2NHKBi1+ey58LG+Mfp8WZv2+z2pAl7hHPSqdzs9BFSu
KVbQ9X7GW9QlZDDM4cKvaa7sM1/VL5vcIATueub2YEPJhgNKgn19M/KicTJoTg0SnIjflhJpNG/q
P7CAp+FXRPlnVrLjQLNwSowk0RTFuTPintX1xlQd0xvSdeWVHqnfdtCQZHA4pefNbo++GO6er68X
JkHaQaf+g4TiaKtgAyG8c0F3RX0wvp1Xv7XrqJrN+g+aTlAdNNFBOmRR2FqO168ut1kjwfYE6/RN
SQPzgSGLIxCvFmylAMcWr5wGj8GBtJByGdcmMl3BVdx87shXqi+07jLZW6/4WdNJTF4/y6UAIuIf
b/DZTFl1ZfKfGufeBAg+Hcwu8WYozny3M2QLMKFsU5ZZYkABKIRW72NKkBFnbbF9pWoLLwbwyqs2
vM5UzHOPuuUDqgF54oEH23LNflE8BSi7aDdUr/dyM1kCwjo6krUlbsoXt+ix0S3b6ZXUa6Ajt1JU
bQ/4U9thXYIe5J2pcfndNFnumiL1ic2wwRfhGirGtzC6JBSxej0V3QfZMhOkDDJtMZ4v8+d9W3V/
bKoxBs364+R9ztHg9eA1pwmhEutz/JXlqdLtyPj0/S+kxMQyYsFc9WopOyYFCECg90o9ZsRlPQKh
WX1mqXZfy4Tx16vdt/RqmdoAkY5ljqG1WmALJKQ6DY+fZ4Z1bTodrGgE03IRm5obC/PbpwXHtlTl
swB9r3cFS12tyPg61TWvLvLP9zREWA50OCkGA8lL9gKmAFCbuPi71EnVegHEENZpsCIVcgED07/7
YWtN8E27XCbL6oFHOtqOecY3xV2ERUKqZPNPAjEP+kcUcyBfBSQIPVAJ206555lWM/+j8HHV08wp
ZdyrqbH/SUt1gTtceArHmIYVT+gKnjvmDHs7DwC3f29QDORwTBAz0WqyUA+2GudLO499kUW4u+eY
hKIadhdKTC6UwGuKioBDlr6kNGbcs7EzWiX/2aTnCH6TZpf6yr16W+ep4Ez/kb2F/ixNg8s/eMtw
lcWH+BbTp/WIoIonr3XPpR4nrjhXyBfaCWYa9jmL633rGfj0vQoK49ne75Tx0+UErnuyG6N9y/39
syi2Gc6/eTpg59Po7QcnqZgY43sD7YW0VgXVGWlPDrmroxfzpnzVZn7ec8qmIrsXV8mVJxMCjwpP
i/8dQm7fvB0lszVev1/YKCvHLJT8ynpk5u4ZrXbLW/LSfkdsclofJDvNhRCDuobuhUmKCLUK0/uz
r5K+GigyRcAYM0BqesAPH3aJ4nNeE3M5FtcBjuUOWOHcwwLnvkwrvpnNhV3djRJ3xgFlFlnGbivL
xgCfR6TRQMIIuX8q5RGBnc4hrYQ6c5vNcv9EDiA9Rh9xQ3JZnMkXNMyOGyYdRsHCmHm8ZmQCknnf
yuTaWEG+cpVjSmbj34gBl1S6KlhxjnnMqkGDGaqyc1Id9oeWVj/dmlUNbkVz3qu4gJms/xeDLQBV
rBXZorYKYjMxfhYCaM0UWG95knBoEOqCfxYVtG58Ek+CerMR2aiA0LO02PrrTJ6VIiIH3WoVfloj
kIFHUPwMy8sGOhO/oQZ6V/6LWy8zvTSn5VZVTYs+MeYuJJ16xkBDTNHvDWYUxsBJ1Q3ux9lxeSPo
y+cMIkp4aGHOXhxbtWx9PJfg478hpin7dTq8ui9bSwRc3tNxBx0AowUR2t8kIrX6QOyhiA9uX5+n
2cda1jD53NehSLrDI4i01PJdJYddDmVy7SCtP+SabUGfR5JC1FZOqBpOQCnNxdekboIHrFCaPaWQ
IBR4TzVlYMgGxIZ/w0B9DrwLxoG1P7cHaNNic/zzFU5X546eeCuD5i6e1vLFiG4q+ZwteT0LAba9
32Jue/AzaWbjPCuErG2hrisx1821wJkuS/tFSKXi8aanJ4jPv3bsIkZenoGzxDpk8Yrf0Rcyw8/5
21lGh9z/gdTQYK1s2AKEXtYFsrg6RiqgGPean8XZbJfDBkPl67F8ObogWGYicyc/0KUnCqFaNyYh
Q94cO52hqhTGSSMbcnqp+lW0tj4aiwmWgVfhQp1Beofi0RqD+IlsdL8b0MJJL8N0iSeEBsXpGxgh
Ozl5b/RrW2UrmHeU624mKySpMxVWgUoP2oUbGMzF8K6feL1hHX1TPWGRH9+2195WPI/aiTV4GvwD
5kubAvIlPJuaB9he9Z/kchf3P/Pg4Ho2ChrIIwj+pog49AFaoJFL7F4ERk5Tcu+7iIlYlCU4p5uV
2/pd1+UhS6kT2Cv9P5bBY2RzAxvTNiC1tPZWZKMRsblo0C1SFtj8PK8KbO35lBUbLU34o83AmT47
UvZqECiE5IwD8RSWYCd0peuVLkYvDCPEyh6HFQTIojfJT1zTfrOwYuwZaqrQEqqQNuMExKi3N373
LjqCuruiXRdze0VY/yWD402wmOKUwKcblqsz46eq063hhQJ6XEXNU6Lg9bYOOVdHBUVu/3X3GRY0
SBad41q+1xvabABOK03Re24KRJkyuG6DyPWIoola96f3T1j7mM2fTJrH1ZG/j4kz6rDsVXhchBb8
V9HmG+z1D82cLdj/D4Ot0jV+FqShbTZO0r4QXC1JcuApJoHDoo2mlVWsv5eHgIatNWztISgERWd4
B7h+VuJ/iXDLJKsvAXHBiBEWZ+8vE4mbipym51HKvgKK8LDyxD4nArUa5Tlf200h2G1v4CQleCTe
XIUYIJmXEZkAHl/+OaYt1vUkSM4vkBEgIvWLelEP3Y+5l2t2kYocJ9lV2+wo6zy8bw1kLtjYWel9
lOYnQtHUJfhTIf8D8ZgNFx20SXmQSp4Iz0gCU6MLHWNt3j/inFhkatpjUOA0X8rtBAKl2Z/nRfC2
N3TGNmFVMejz8zPAccypdH2HOg1RtXAoSRtQFiY+++mIO4sCOydxWF8IuKWEd2H9ZVGWF9NoGTy6
646tGQ1vXqLLMVWlQwe/+WaX71J55RUgpcYBggI8Av2+GstEqkNQ4yHpUVOa6pMJCSjQ9eqCdBhQ
V0sFpFgA6HsPKRBL2cQLyxjn/tbEsPIBw08sF+Uuilb2gsatmb37p02QAmh4qB2QJb9lq2WX6j5g
GVo9TIiS5+m6yWyqVN98Z7pCYAM+r/AZWXeS9sU1/nJRrsFuzsgEQ+tLdAwh2CKb1IxWhoBQ24Sb
n+Ge+c15QbKjc5elGGjrCkztj0aCEFzOpOabmGT5acuFZizOIYhkyGnHL3tERsDMnK6rohz8YEgN
doJzOK0iRta2oJFUgiPJdJfkkv5n4T0vJrhL02tZbTAfxxhCVuBy6L5R+LyQlIPnKU+/E/d7SLCw
Fz3OfQDUJok/FTx8J8SyOFLLXpXKpcuLXCLaoAVei3KumCY2BtY0F2YZYFwIBHlGLlDC2CCK17s9
0gkW0JEsd4sGF/8Vm0w9vhw8kkNEwWtijz44n2DArAZ7i/jeo3jMk1hivvq8LFZGxJEBPbfuw3go
rE6fGIaQNG1Kq+GgxCe7uQq7dGiKjqrVEx8KE19JBfIPnPV5F2gch5sssMsn1qQEygeTG9eqA832
V43NJK29SVHGxJ859cHlsFJS8q5P1dKpcjZ3JxL1zvyjzdrFr54SNVQOWj0bNedhDukfSj7YCnXe
sO8BXxupXIAsAO8pKyO9gehZJmLoSq4uImIhLdFu4r8ExUfoIrvD2OkgWaSOcXgAax7BM63Q22RA
EGa4lNGW5PxtUFuV537w1i6svItFuYSv7ZO6L0fyK1Z7hNXOL7fG4EYfA/pE/XmruK72/rVJODj7
a3sJI/Jw90dD2EVpxLTcQhdlqbHES2lVabhIiTfaYJqhLWh2UI2Df0lO2/6Ra3r4CdwV5Clqc0Up
vI5xxzL3P5kgYRrUTJLb37W0EDwOniuCWyWtl/BuGz0Jz4KtX9EVMLBF3/p+eUnSGOt+WGAVz+aZ
Y6XmTKCZ5qJVABF7EDPpBZWC3pxZAtto2VBK4nU4rW4VH9t+wznU1aZqAvYsKK9z6WbROvuPBPn+
O2gMG6IJiP/wAnsrYhSkdtFlvy3W+Oar9ebw96njZlmK5E6KLcunfTLmhoToEms+eB+77zzXgdJt
smpJN1PYkhcsrVP5arEftEYZbeb1oxZK+xMlZUBhRc2/vG4zy2l4lZxnDxX6DsK/nbHFx1FkYyEl
U3IlqvPkUXJIMp6x3MWFjwXs6/Mvlc2EpNFKruD8l+mfRs6Kwi0oKfv+ZoYIM30BrENcNXTQ2D5m
77aVz+kPeRxa+USFxW6HGwLi0PTESfVlzDo0jnnfif7IdaD+pP7+MrZOxMZQ2BuI31uCatWBgaac
SeIkb0EiqU1zURAWf3KODCJ0hwpfoYFHFnhSp0jb9tdNYvI1O6PUAgMvQDnHhfOtnh96Iq8p0DtD
K5BpeDsocpMvqo0P0RszeYYfsUw9RIeMivTwxPbeL+cVIFVyou/iDTYxmY2flwt9VpEgpPW12XHk
ixQcWzOf/2ghvnjmFn+Fh74Avc1ElUUMNRFPXlgVzTIy2j7NBxn68mOLq/WEfrl+jY1HLadJXg7D
KG4rdNxSQ+UnlQLsOWILmi3d6XAJ7nNhekfve4fS3/YS5ezZ6YE3UlFSowm0V5gQxA/M0xCRY096
wZBYl73kb3WMNK1Uf+lGlv549XKIWM6xp0RbU1U3k0rqRHil+fha8qW/u6nS79jRusD923Puj+zB
ew7UGh8Wiu4XCEcoqeS8eh5B4NUzas6gqRQF+ltlSipvUqv38sH/3ycdgMvnif8JDUMxLSDFrB6R
InTnA9qALznV3HBXVuWrGLpsdVPb2bLARhBkmS3W/jHq18r/bUL6LCH0VHn/k1vmpzEIGpuq6KQZ
n3G5KDQzX4WiUU0knXdpFWbCn3dEBTJ8eNJtGaTwy6t5nUyQy4CcJBqAgGGATSUVhspVJ+w7pkgA
zMzRQARuO/Ae32TxRSrsHd/dRr17L6cIhoVXPg8+WU2LTXm2ECHM6OaGPwfDmmfX13u0rS8V6az+
AoIzL4uUGX5XYsjHGHz9eIt5OqOk0/EhFIy4QFPgM8PSvIR6URXX4Z9RMGzeiT3jDeqcTkLICMat
9RblSsTU7zwxDDC1jBP018EeDZRY+eJYYFTH/gGFbkCPZ6HbphhIH2V/ZoBWPJor9tY0N90pnumc
qc0vB8LjzSl+XH3gZeWUrzCDLFTNYIaz2jpbmUeJw3RNpzjJmBmJSzIT09aRcXeDzH/7ktWD9eq+
bkukVg/T8w4boMSIj5h0k9J31JoJatoPY48QFuzOl2WguRa73JmwZ2A0yhjagP67jDxjXzIKKaNP
SkSkQ4hiISnPYN2UvQuLStpCdx7zA7t0QlpJkcE+6Kr6UkZCsGpWwQJqFIrh+MIfUL9YZpzEuSOA
fOhAgiV0xpodZ7ttc9KOzl4XQwp9zj5y+5KKx+4YhZgXSGqt5rM14vH7tJlSPWgT5doe8xezXIeX
kdl3q1BasK5krM/P2cglpgUa/NVbAxqHMDyhMuNIYjhGmIn2MTAiRZeaOC6XE0DGGso1kVCjHB3E
TTGYpfiAUPIlWe6MtMx6MOjrkYoNhiirgnUEoo6GxxcaBeEl3TR50I+Rt/7PIlG0zNbdnTBwZky7
SaS/1lF7wDT8JV9dy4DHtFv003AV+id/+Ynupb8k2G+LZX9UL4VfmDD7rNUcI9TOxOTVfgafN+ol
yLfJQJxSva0Bih9Z8sLDOFyzilICEyEE39bdmsqCo6+YMDaYwD3QEsgSVgNmb/VWlmGk1rOMmHKl
IRQqbe4X3BIO5OHXRQ5yyUO1QBCG3ExdMfRwSTYeK6QM6lmtbeZyGkPB3iq93RCzW/gBfcA60u5H
poIMYyPE2/7nMOKybJ/GItMFBcpxrdXDWUQ+RRNuhMZHGPSWrgGKozfekDvJxcYag12geJLO3TI9
gr5jZgRgmVdHaZnePqeyBU6aCg39U0/IASmLCxe4Bd+U+QF6Q5QDoS6ASGkSrjohZP9Zr/8lQCGK
wHnjlNrb0evRZTof9u6id1pi2oFWVwEObU+WjxiBravUL4Xy+7h/vFb3vZnpJJcTWFQH75+9mWDC
Y4UaJXYyJwSwfxvFhwryuqT3I304xfclN9eW7COzWnljJ8E/Ch7SFEAgpptZUWuysUkOqJ4iYAky
dGGLmarNUegirV1bt4H0B30ahcbm5bgGmXGGt6vpKyk+O3YsZHdLxzI5u3fT0ShZtN4i1w3FOMdL
yWdoNQS/AdaeiLH1Pc2L88pwhGOd1TnTKvwIXUZU/WOns7BKF7fkHI55NHXakDOhMl4lrHoFucug
EjpeNMaP0OPl75CPChw2aEVZWWkLSMlVTbPn3FgJmTpV+fyIarxPGS7bX5uZYuawwNETnlY+FDk+
XS2l9nQKc9Qgx2boEHljlBp4yEjZq6FlRdEKH71OKT1osf7qHejruZfdnmpcuyQ18p76U/m/IGB/
uHTMNuIBs3CoQGKFf8mjqucz8NZMZv8uT6TX/5MKen7d2Pd5esiXHhIcXqiXnvmMp8en6XbFGbc/
bmkeW8LizVy+h6mfN/yRJtJM7gfFJmM7hpZhYvchbNFFJORowI3PCM0cjURQL9kjDFsnwD/RNAqC
0e5tlqtDOaRzK1VOpVJGfNjn3BuRdMKb2yCmNIyG5hIJWo05MnJim7uYtk+5TsFCHuxDOaDaAEoE
aCYIv2Bie0Ei6WCPqcr1IrjFZkaUV4bBqwTlN10tbSP3xGZ22X+uhhm/LUaoongdmxGtN39GiFFg
y/Z3Jc3jpVx+QnVmig1lMfmdMXTs7g1rf6JXx1BhSuwBxBXZvy7535taL+55N8241ALqaDPA87/5
DZYxBqK+umjc1Bu6avmNZjIajzTMi+/96fvnGIydPtzHYqj0Mbru0WetlyJ9/hluHZXC4j8kD3w+
GiZV8OFPblrE03A8qqQrhKtUf/PLuhwJ1T67Us4IcFzNmVQzpf1u54JCWRzrA/YbwMIE3fg57aH+
NFDYE4vDSu9xJf/3lHPtQzGdUR3bIxsZatH/Rt5LuWqDjv4WQOTvMNV8yqXqq8RxeePJW7n+vY9G
fD2/YC4IC3xVdu2YjGyVGI62c77qiLQ4Ntr6jW9xo1NsDo5TyfPWBffkNdD0RzJuZfDYA1iWNvkC
sQTYm/1SCoY1M/JKYfdoBnfxcsXdrqXA+QL8uOnJE5TSe/sdN9OZVbMNU0eNEkYdySb0S0nDu0Cn
IQV/fw2//iVhvrrMyvjQcBVMA2RTklynCRebL1XOBlugsxH2FuaOrdX2p4lcnS8e/YDxxPITmML4
2pxxnXhUrpiuU3gEdzBwFDiRgbmvVb7Qj3hhsQC30G0KvstGgPzQKEoUxGfpxEgnYPlYb3MfEGmw
CZJv3duJTjJ+OagLp4X12W1X1SvR5QgyKdBGx9oDgUgpmff5ph/hD2EIDQ/45ttfZDq6RsyqNFVH
Hz7cstY7u5+4kXR48QBhxiH0SyAmsX3/jy/jimlGpPCnvP78lTPwAd10MOqksEi1zl6ob4/mhoej
bN9gN6Jd4ycjrYKe7OrzC7wOVTkGYUnGuSWgB/rHO9au766BfdlASO0DgZXx7Y7HnNGdnA8uDtKJ
tiJherAsYKcZn0ke06xSOQt33FLKsMYXQHKehvzdAgWdQz+yo0uM8JmiNCGjtVqLTAYW1/Sk2zYu
phuvM7Iupfmxi+dClNuqc5Qii6S2kkFXPF/Tl9adVugBQHBYldhvqEWiHsszH5X/1oI+jlyG/p2o
ZgQclaxSRuCH4tA5POYCRx47pAtR+i1i7t63hquIzD4S/vk5yjTlLrmN5g5xeKC9HVyZU2XYZfEW
xqhbbnJCuVRfVE874KN5l06CH+ruG1c0H/J/5jo4ltAKIRlxTkcDyBTVED1KvrFvZkC9M0r3cjtz
uVt9Hyk4eYLOzE+vps+m0JRDTOC6Q4P8zLuH4XqhiZqqbni7d3GPldyDcKRnsTwkZiLU/ErqfKVf
59NSJK388b0H69EAhJXgvjgc+JWRo1gUXo+I21CsHJsQtQGbuZD1EBASpbFzJjRn2Uj5CNmQcyfq
BDBwM3E9mLFsR3Dn56jidTLyXMD4oVeJAyNzpOW+F9XCjFlu64YIwEQX2NYNOduYehqJtIKUrHVO
ot5mo7SZPCWFOS5cpdv0QFceTN6jug9zYaAPSiSt8E0UcO3YWmPz2rnknTjnukYimAX2r5hb2tr7
dnpUtG4jiPQlYCN5wVU57L6Y4eb8685Avu/W9EYcNh9y0gazXacdcOOQNEXTBs6nsyR25UKCFTdR
BL5wpg8xxDgaiE1l6ODXwSZyAoXB2kDjaOpX3uXOgI86/IK25YikbFTT4Jj5HiO4jI/ST4vrncqd
D/8xGovzdSAtXZIARPe81RrGlRbYc0FZobDHoYgNO6VXrhwepB/M8xKd25cUNGWGT/HFk6bNe7Zh
hFc11zpOsyJqwCJfA3l7n5xGvMXmJNRWKTz6LciOTgH8WNbxDNuEjAkhWrfOEQcEIvACvmtdfvzO
E4LANx/B1/8B+VCqaps3DIRlqeSf3sJFkpvvtfWlbdS8BcAsOz9cwWeenR1oOmapuODbludJjXyH
i61O6xGCyZKuLoBhUTxQdwXjFdje9xUjkYJPG79Ye5iLvzRZRW/EQds6gutT7RtGqKRPaNMLBzTs
07XAO4Q9p3HxSRgLKs/ghdjTw2DnBaKTmtQeSU2u/kLuj9IozV84DzTAI6MtGmSaiaxjJ0+244XD
aA/0W6NdtlrLCM9cKE3rmueCfN3CKbCu93SFysh2FEZwQJ8VARoYlMPkZnJqVUFgtQ55AxdnmyYq
uKybxVIH66YyJSgYdG2cSl1i1Kv9B1lDisEJxhaoVSgrXo5iT4OhMStRVKEsdotScr7hA/+QYHD1
B8QXUvNPQ5E+CO3RGDCzTmzmn/P4J71QhT43mju0ievtrExQJ0fmMpkNew3VXJ060s9t2cMd1Yb7
m7mUtkYutljmyXgjRQVmpUXNFKle2tr3Uc1VfZhqUTQbkuCwCUYg5begDGf6dk+C4R9D1RmgmEQD
VTpibMUneNxc/Rr5CF0YjzLZoVPR0e24Olv7yiJNrhk2a8TE0OGg2ywwv5D8EBKHgnl+q6D002Hs
F8S1KMcalmwLCk2k/tw8HPjz5MOtZusKvHtymLycEdrkwvcBlJz7GBe3kHccj1n/cHK/xRiaxktD
/t78sgzR845tMc2KYcFOmaTWfcdPPazasAJ+r9WcxnO09Wn1/zt64psfUyfmOSxNuU11ejo7YV+A
PKG90T4QH7JnSbGI8YRprBCIZKkr9VZ2WjRVlVoohLzW4vtdp5k6RQOUirCFPl+egj+XIe8LMLAL
k8yHt+OURgGuHgxKJ+ikoL7y+o1unJLX8iUmQV4P/yYWX6V+H+hHVEW1BR5Flz3ByjtRjHPEFyHL
jFQk6jcdc2Yts7KVH3Bd/H06R4eGQo2XzFTPAwY6BQ0NmqLSDdeCHL9ohc+S12d69dhCfgrrPfeo
qwS/jin3wbyXRfpfS+xtI4xMsKJV58C2/4xtyBepLKz2ayo56b/SO06JNSz7orkqIzs88TUUH3S3
ZRCut0O/oLUt7mZltK2TiMeubOJLy9yMdYaRE6AMj98xh8Zhcvw6UVcPml2KmnqA73ImrsfHXlLZ
359IDBuy6IE5bgZ4T8kdXUdyL31O+/lcsbV9MD9/wXWtV1WeM6vsQVK9XxfZT9L72KAaryFSywGu
LWMqT4o+N9t4j1pB23nW9AkheiN83frxFqb4XYeXxCIe+lVu9IodJUVIyEs7eAbYzNJGf/c7EhyT
pRUXCXrFNvflypMHX3pj5NN/E9O/wj7iKrsjg1HFyT2plhIAjLgDTU96JnVVGvm9/Sosm0rW1AgD
39RIv+RPn3ZwXcZLDyecMlcHNiIl0Skoa99zLrHLmeeCf+4DtKBMCxQVz0j/G1/qi74b31GIvDgp
lD1gsh2k6qUUQqx3IepSEzofZuQxqJ403Vd0EVJOrjIWd60rKuuUSb9Pt8bGCXzb9mLBu9zyAAiz
TnHEbQnl4UXqy45xYTbr4FptJLpA1UAton3S1VRaZm5D6D5RC4F+u1n02o6L8DW2UwJVOr30QaWQ
Rq2epiKqY6nZYDcorgAYO/vJRtJYMJjFrN03By8FUhyQX20/GcMURBywt3T/QB3ijFOqK7ghLb62
52D0aFkTpqil6qWS75w+PIIKOU1ogUV5S1YuvY/sZM9f4PegstDeY0UIcFchJhWcG46Bp5OsZBoH
Hj1ebpTTZJemmWQtabAgpNmujwexQLFsotSBRi+ga9bDC5hng3heqZgyhWOlY/jpMhgFex5lLSif
00VXuci4ytNH94/2JPbQfFeCEUcFqL/GeMnVH3omeyQHiFliodlAMvkQLizAP9w4lLnk8gr+X6AH
eOmsoJG81px2tNjJ/SLM0ygSch6cidHL/mHQsKbBSRZYGSFSsXZEbyhtq3rgW5LsX0B9zySdRHPW
2EOMulQVQRepmCq8Gl2hOBuKjjRHIETQm8rjWbhpUwHMi9fu0BaoGa+zDP5/SuAUcpFqPffayPp3
YPSnpsQdmWUgxuEBPd84RU1esIjY5Oxk0ZqitwR/vLRdUeXJJqnMqdGvg/152cqcIxkXJhJyb8Pp
HCm6/zCFnS/ATBjjXyEu6LTujDvt/AzcOUK28OHFCziDUehIC2h00F41hJyu0d/aGQAvBmA6F0bd
sT3gBi1IykUk6TaVj8Xyf8M9peLV//Xtu4MsjlkdYamjDcUgAUozn+OpjGkSaO6ut7OzabHsD4Bj
9J2BbAlF/+w4OTagD2cR8LFEFHC7kNzTQtXa1SuKo+yr0NfPV91GqiIa2szlAfGQXn90Z+baIbce
Eyrcz0XWHQgK1eL4E7opFxapSZtdKlWoEBC0yAyvv+vPSeHgPalgBS15Wiu4hSlPa9I+A2y9M7eR
W593NEg8gFwO75cqr3CCRH899ZTEk/suvofIwWUhsWVAQwmGrKmIv4zVwgA4vS1OXDTjgohSbrZK
psqoRd7Uy80P3bINcH82tdNW2Vht8LkBE11JPfwPKObcQ9/UB0jcueXBCEQ+rg9GGKGZPPJDJVNh
lsx7h8Idxs7hsMGW3jdLHmTzfOWAi2lQ49XT6TLxiRMnkqMla3oe4Omvl1jdVoMNFwDo3Ov/VVB3
dDY9iCIyYPiDJITX8NTiDX3UGYXL5bhLVXu4rizR883yPRUGQ2hNg2/k4E/AxmJeucxij9DQ9q8v
dl+0tXFJ7UBI6qpyBFPFrhk9xviNeKVW46N/BEyla+v99JPBvbL8b0SnWiasR3If6NLESTUG47Np
184YuESpWdfh8fiCJChMtV3J9p2CayPHv6vY0Noy3PaDr2EuNyl5zFAY1c2RKtkbc1s/+zzs0mGx
izcGcn81QiiAebCyiCOOZTNQHqBOrJtKwG5peSU8mVTswTZ4uIK91w6a72lzSfg6EWySZfFqxnKE
KMSCyEIhTzXsebdWrffPSrMENK5E6RW7DDNh/roSd+SvCve2dlX1z5rhirlJtXHmBnqDQjBfHFvx
ldTQt/6TjzCOidknWY8Ur/RdexB405TbRDmssxRNQiC0DMoA1ES7WVRJEwVnYuY2csU/fFhuxlv6
q5rXWJKUTin0c+XjNiXdyubUY9Ks26cliSaZffQ8mebrv58XHH2+4esSxtdEES10eJepC9TBGouM
SDfdQ3tIyxikFERXbfg2PBC12EqLgvj9DCPkkJaRPbZzlNZoMVuebRSuVrQ1bcQU4tlK6iv+Nb02
ChYnC0VJasXZ4Qtnas1j3AkZD/bXEGMzQwLfD2wvo7njp7fWWNmTUARy3bkO1j+P9XKOrRDcH+EE
Mf0Ls2tScn6pj1sj2kt8MPJuxQeRKnaRTpMYioaprUWmBVELIdYuVuj9w0ZfQJeL1d8bx5871MnT
mBDZlkvLBsyQkCmg+9jzpBC4dS/yBKOxSp1j/DW7CQyegNNzwGM/dbA5or6bmIwmNCnWwqoNeIpV
eFyEHDxy7gwcybMfyQ6h0/41xpGtp4utR3R9YZkhE1UoAKajkRr/hsYKASZIsBg1ayx67hHdDxme
PzNgv/JyGY8B/7/iXuIqSYi6qyTV5/GApvkceFEtoRb4//TuJBJA1Y+FovP2sTOx3v6FvFL5CAVb
Ne9PirGAuj9aGsV/SfYCwNFrvcjmMVmbW0pkS1bFO3msg93SOSeWMWCEGrsI6DrKJtXlxOaJSdja
o0cHN68l0DtmEQbCuQcl9EpGhIO1KrBuZtFIvGIjGtw9mJ4Dplhfore+eZrEDvO6q80joLBF6g8N
PEJNRJwYctBIw5dDeVJQDPKJKqlOzawVO7mMBS+PftAc3kRctNH48AOYZZcEanZpQQ+y+5/rrXXZ
X6PVfs1VCgHJvzxEoOD7FE2oomTuRrNlZ0eldFYcWVsa9YP84AFE8MdBdZghSJ48/n70QHrKXZVq
mRD9KDVEik4VvTJzqChhsnDwvqHtXJ5jLC0wanyFQXZE8qcyNsv+FqW5jr4tw8cceIC2Z2rw0F8C
tCs5F33xyZDELA14WEQB89XbErAmNCH+kriE4tLQIKSgOAx2CVyGVqQ9bAjcSVWHkcEwyCy+7h7a
IvH9JdhhdCgBslIHfh+6FwQqBhBrqA2JtgfgIauIn+iGt2krjrWPkoz28UoQMHE0e0WA1m5DLWqR
twXQKvgGqiN+RKedscGq/4Dl4nc/g50eoVNsNFqsljSFyZPgF6zR1NVy1/SOgQPMrpaYwpyY+hLe
LDBOZIrf72okHBd+mSQnO9DAJXiG3Gxq9FHCgFPJSuLb1jKIWa3x1YPhKzddIIdB5K+fOfOHoMbI
JSLJvCM+Ek0xgEf26DshOhtwIdgTG8RE34mspJvC/bjuVzhyBXiKGjGHusXwRxH6E+RmWFq6bq1j
XvXLBfiCL/kiDuwSm9p76jvBScYqNbOvn5FUVSBLgFWCMKYPZ01rQHZLaYJDgx9z8b1FOBI/t/yn
KutCjdpvZLcathaYWqF5wN/Y0uR4U49YAyh33rdf7st4evbOMw7YWakPQbgZ77QbnCt0Khy+cjsU
wCe5Rh+nvuzGEw8kVrKerBVSRk+ZS93qVZRUBRGm+828cT0R37iMa4Ly6DhwrB0GuICR8nbSKNMM
b1TcbuYww7LOpOIMa/3bLLDOII8WJihoTuQxarCeVXAVtMjmYPHARAKHHZHBfFWKth/8gXhrHlsI
Blg5Zs176pIfXE2BK0ZHjtgvxCAOTZAVC7NmI2D3wU5ak6IlTiMf1ceSJSjo0Dy6TTiDcXjhzZ6T
zLiha3GcRLNr3F20SC7MEo3BI5aMU54jdODiiTuwo2B6w+E18KbYiOgCll78eS5AaX0WjdwyHDXm
tRkLR7RND1PjiFu0eCTWtqXmSGvbvPwEVEmWQlz9H6E6esjvMTbBw49MORkeyU+8F01as/yv9bxS
wXXawTtKbwuAPu9QuSR/bNM7jOpg83RP73YEKktso1dReGqA3DT9EZ1pyZKU7S+IH2JZuYp7sT3y
EeNKAOYr5QHP5nvcgzMRE5Ydax45rggOi1Z5BFElNn5QwFrV0WWHhJSN+3nMLxHjKLrcwcmhbnl0
BrII3WWiHJf8oGKL16S1n8qLFU05YU6wlkt1MIJqwSgawbPlaTjiJzIzAEHD22hcfrLJf1GNwaoC
YZxD5uvMQ2zbTr8P/ta0WtQ8JVY7fJK1cIUm2OqTniambYiBuVIRfWSyjKehIHYwS0mU3V6hp9L2
DRwc/0P/Mh/m3/PMFMpqsCbCqMM4Oe/dALU5X9n8uC906kLks+oofoRy7V6habem7oIMVG29/tqA
m4RWcDSyIutKbWEutAxkP2nygQ1AEMLlp2UU32Lqta5LV3rw7LtrOgMpfTtAknt1N0Rjnu6K4twY
0n861qiMTJ7+R9n09CBv+5yPOSsiJ/ZVyaB1LISXqeW+JygFbyw9qD+5pyEo9RMj06nd11s6GFI7
RnQI+WM4PpWyQLZktMlApr6r58a/rFln1MgPizJN0qAFtDDQgxMNJoOjRKPefLydeLGL/3UEebkw
o7bfT+EWsNHtP8hw93aEXus4fjDN6riQs3GgYERPp05HzdziuWD48PZbyVCRNvxrOQUlC6YJhTAD
Ic20la0o530dcKnosAiDd2djfqnN3F40WUWAKMV13+ILlBRJCYOjxSA6M/zikmQrK2zmijSiahsD
4j781Fvxd2iMtwpsPsD/YF5kcR9H/mnqeKAAxdLVfafOnKi2tJDxU9/d2huKOim/AkSGUy0BWF46
hLaJGv3104iwyVl1zqlx+s4lTFgkyOFqIDUT4Skl3xez9FHV7ooABGIgb2hOB113lYvZY4Q/ZztN
9Qj0bwDuAdWNtr7hV+X6BejSC0q1eZb7ABBdIM+hRDtpzPiKqD/9cNFPNBeLtJqZTtGSR3lqVjDo
vR58N7tZ5SV5Ls/hl/uWPewWTNgwOptZGehc6oiqnWm+xY6FglgaVBHi2x+lUe51xJ3OnyyaXE4p
q6X9ywS5VIJ4s4juflM4F5o/RGEx3zRkL5iYIXD6Sg1QoG2MKSgXnLizd1fIehRUaeK4TYm3pAPh
o30qu/oRis9GJVSh0/jlvNDWtGNiAmB1V1i+fLXtPTPIxQKpLAoRNvbKfyxJGCWuEqTBnGZAefI2
sZAY6AdZi44/eOf6MRM93frcdO9bzl/PAwUgmu5SHYxHA8B0GMisAVVKRHRbUogMGjo8pT5/YYeV
jdOQ9rFPcogPYHnUvahmXd6tYBJOvlJZTmesxCkSnbKWbcUBnDax2ALipiOz2ExmkUEaCl7QM9RS
zmHYd3jJM9AJ56QeQmuuDMSeqqxe+uo7ktBEmhohUNpA5UFBHdHKNcR391nyps0xOH1J2jVJ5f7A
DeI4OwLHfAS4LvXVOdMNPLlAFFXNVVVxMTkgcR5gWnWyLhZyi28BxNsdKhpJQjjLF32UcIZrfweT
dZGiRCbItNVW8fQ16V+Ceh1fIUIYTv5B99IU8fXW6ZeCSuwsLzcQpnve4AZv1iHbQwIo23ydN7gW
szSxiYbDvtZZs07Wmbf2nNtcnsH0ZUP6zRSQ23LgW7oRzB2wYJIExHfHHLTrmQ9arrQgZ27vt+zZ
BuIIvXQQoguovZD/QcCH6fKqsLBVmhHgx25Cfy1K5DEdOH3jImpnD6onTzHkPO2cSwgoX9CN5Y6Q
Px62BLYk7yjM9Gny0Joquc7VBe1Xk6O1mdrHdyLIpPKbUH6sMC8EhEpseE65FCuJTUwHXAKdjYhI
+LoVxo7WrUsdOS6HgyPdk77IiI6TN6nNodb8u5pRHIGs9bOS3YGSAXKpb58jd7G3b5I016jANTwn
mUztaReJB+rYeE5u8OlOKSqk9VQl8Xp6UBka3vGKJW/WupuXCBIydBFiqhL++rVLDl76jQAXS9Kc
RIbqiXouNKbqVfNMSO4N5MI39ozzVIJfOPamIX4/e2uySdrp9KVSLorr9qQm+K+5usM6y8vrzq5S
qC0erH2vvmD3RcBBrp4jBoD3SlLYzf9iINCgukCkL7NC2TaYYoOyI/lfZ27ZCK2XLHM1dqEhV2mb
3PgAO9PYwBoqYPsUigcQjbo/kFt7JKBTsJAloWK5WiswXKL6r5wJrjH1rb37OuhcoWMrk819LjWN
JAvJx1yLl/0cMEt4OwUqoOdGZUl+RaZFJ68+hUPDCKDsYjJL0v8UbY80SZhqBEDWwetHvVWIs0YT
HkmwYJD1mYOSNrC3zbHWqkKuPHAa1CiAuItwL4jtIb8qJIXfrQe0hNLXgS1s50ydtOF3xVBSPLDa
wFygjXlLCH9GkRlJho4MNYzI1ny6TlhuQx9+4GqCbRJVS7/+DaoagU1IfSnnoKViIO4qYjkKkdya
UWYQc1vfGjCDd7nd2Rs3NRdYc4e1kKerp+l73/AWgfN5lSHZuLTr3eeyv7lhTO9IWD2tXORMfuyL
nobcDi3JLG0DG+U8wBsU7ShvM5RWpJ++ig/6h+6rHKrZf1Oxv9519Tiy82St4Mg52BGqTyWqrtly
uh+eV4d1M3hYysDn0JMgeu7ASahtL7QMK+l1FURwc8JgFAShub9rAeN/xP2KzG+GLsoTu7SWj7oV
GPCLdt/zttDFae9+MDEHQ3SGyakUOPcoUwQaWiPX8sbLLnXN92MSufZxZVoyfoFQXVESU7j/RI4q
KVbVk6+F/8NG4dMLxMdEeF4WjsyhyNtGATLH99v8vtmvB7A1C+cYDXOPHSfv0kE2joZLzMmt7nnd
+4qeXdZ/8p017UIVaWj7F8H9dxQwD+HhNLDlq5znUfepAr7bZed3UqzYy36Ipbq7dkcA+aeMg/Pg
VsIl1MXreX2XJujaZoZQbINFAFYAQ5Cnzt3fYblDQOeC1St/VowU5xOdb/8DaQyGiuHBUdx1UKGr
93tNadJ5aT60uepiVVfeyWv0sFs5NJg//tIavIzr9VKe/4vkzA7X7jrBgIykmyy6z29/QAwI+hRC
us2nlGksDAMLDcLAK+FTCGyMlu9m9NsF11VyDtUiUzrWquescgmtxTm2ucUvxcPg6q8h/VIP/vNI
oj0n9C2EgsxnrXooi7D4oUmGdA+73TDFDgHkpjeGYYYNlEHHFfjwWFfDt2U/o7d4FhYiPiPCNIRs
HhJD/ZFq3jSFW1DX41SR5fHTppkNCP9eHMcRdSwAvPt59XTlq6/HzZ9SrSQcDG8atrCtIsQ+epcg
BpwZUsBkphA3ho+qz3EaT+vflr6PovEF/4NYhukJ5pdz0RsvQPOxb2yExCfI0hCUkxrapntq+Xua
EQVukjWcoUkLDKnqliEmAmUDAGiDM3R8p3rwBgbNie9859A2VJsTh7QV3MwoEBUBaGlYZ1QrSGtX
AN+aNnrGLjCksHNsWEE8A59I803qZHVXiQxUrGGrxu8beWH8XVpnN3N71Jh+wtxR4LgM6SCwh1E3
62D0RACnwkPrBqYVULc5yJML0bERTVaE+LNU3xzO9C217J+AS836RCSkaZNapOiLujfDP4i4sH1p
H6Jj+ju+igvdlmhkn0SZjtJzQyhLM5VbzFJ/vSnE4mYr86zRBUA9ro1Ig/drTmPNWJ0jvRwPQniv
SWedsRek6S7MT3aoWyY990rajIp16FU6sW3tICB6pHg33jj/IQZEWBlHoqBII6MNLkt224IYdVnK
z9jrCoinBwAeQ3M71j5C5JdNd1DcNRJmQHE6NrI2bnJBCx9snIlUfCv2t8Fl7Es6LlUI+Ev4fTvY
iXnOXCKWENiJ/3Rq2zP2tsqAvSzqOqkjG7B33FoCiYT+EPjLaobS1RJKPKf3xKcJuxtDeKD/rZqx
jIax2lUne88ksE1uzd+VJkjnNBFA5Ep7E0uoGTXpeTcW31bTg6NhpCT0YyuEbeJdreIdaV+lLZNE
gaGj2flupVo/SiwdSm41ms3daWUQNTtH81svM+nxNCCR3mmZa7Fx3trYGX1sJ2S00PhW00TzXggV
2vRWSziUGc4YGUvJlJaFat8IQWDbncjcwKL48XO9iumNJnbgXpicqAlQfm3nooLIb9uYlktB6teM
ymP7DiqrmdG9UQv3JWW95yH81enJBydfnjkocUo/wS615mthNblS6bYbrQaGc2T9p+MMQnezYFQz
AkIXUodzchXmocEWOiBJrA6p4V9TvB6jWfrpHO6GDimJLV1kvGjUoO9+OmbIMhRdBsVcoO2HCK93
hPFt9aWRBiT5ShyqLqnh99YjAVNn140nYZQX35Ite4naxcH8pzL+/Ra3yNZ9HefwG15kzAY3lJHm
LtV/W0LQ38nP3Rk/A4uAESmC09rck8QHbdtXERI8T0UGkl3sO6wOGq7D1dUXVETVi9PCXdSVc9H5
RP5RdIdfDnGWHzjZ7yFTADcESDS07twjSUVsAaLV55mkNa+KmcWFZyrpxi4q3O6pEvJaYx0ItbF3
Rr4CoHMb7MJkjCIH6NnP8XSaKL1dPJi8y+Ih0BRV6ZLzqaPmXKGvU5Az1pm7WJsM7Lh5AdCkJEgz
Sca/jRb9RhbhjQX7F82CWIqDNuvixbL4KeKMJagDEMG/PjH2p4eGrI9QVWuw/NazV3tYhQhXj/4f
LS6BjLPCiqVMg+mt2UgOJN/ZFL21qQhKU3i19E5zZrWnZ7gf7EPM3hiYWAEAN2cYXItqxtOoFFO2
gohAHj3H6sozGPpION+570rdGJApQiElEDLGOKG2L4US0EsQwNVf4+6c/6b6veB0oapknVSLYHu8
1RmdrN5tXBiTDsO1Ezz8oZKfHlhlc3o5O6e5j4QaYJDOWVoZYsfhbFHbgdw4h+I27Azxfm7RNyOP
D43l89eMnvW7+9zFfofc+WUZivLK/2aIgNXEOi7ov14auN1QR4m03qDFSe8icK1ic+HLw/9EBnyD
u4QclfF3zs/ai2e29JfJdjnndgvrLCUOPsG1ggzVeSVlhvkF6+B7DdJQvepGndUkKT/LJ2CqBJex
3amUL0AR7uIsjvGixXKIKjK6B4ZNqLPB6wYmuO9UbVB9hiK8RXBdz3RTjEpCiOZW+BZMQ0prPjuU
+KVCO5EuLCNkI1ya1DdJnccuVivXNnV6M2/0bAqi59WI+I2AyTd5ERh5WyfX6PcMEM+UPYqFB7KZ
YI9j4S9IgKns6gnabon3gKDvUYx+VxbSMURWJkGdoMKuoVt8buMUNAi3/WEGEDfWCcWB7NI4StuV
J3nRAciSlZGYD0Uz5bM+xh+jcwCdf8RSrugsJ+YTiTx4GfEhA429EouWbyHzWEzGHBeq21roCprM
biz9TcwErlqCWGeNf5WLI6+MJH7osOZCfY1dR7IErgtgit225y0ey48sBL/Uko6N3mWkzp5GHrxJ
EUewxqb0Vw3gevrPUiarU+Da2lDrUb8xy8Xy2vxQLr0hoKBARWoQQfXRVkbO+Ehih0drV8UBB3r6
yg4jVrIzGi7ZDxfyha6wQabLSSUxAQwVFxX8aRTT51dc02QPVR4hhh/covGmSQCAANUJeiBvh3qy
RWnUvT6dXvfLGwQ2R67cZk0AywpkQXJxR4gCD7KlBkwNZjWmAuS5JCbm/3ehEtVKRXho3yYcJ4fN
Mr8iCa4nOpAV0mc/x/txmUWIhxBvhGDq5Bviyx8qbsrczGIOwMZTiPMHkhz62ULvPJnlpOl0zLHL
D3YYUYP+guMGNT2KrMgkf7WyTXiadCq6iexMP+DAF4SR6o+4m0qxAb9Io4ORzgrDX4Y0mQNStC1d
GTH9xKRKavgA8rMQHPIuXRmiFFgUv5es1Sf11I6njhMYhw/jgBbdrNJbSDQOJBW+VrbS5+XNChGl
rVewSp2xN+9WpN25JuXy4whKYCW9zCHZiMdr3n4T+/SXlpW6nUoc9R/8JwjzFIozK7C9ETlDIsAR
2aVo/isKED7YlrJhJaWqKF8da3VDUYaOvFfDffhcHUnWo90jzZ0lDbxRJrjeZ9nFBphEB8syqkbM
3iMRrhoMc5D6UREScSEmdsG2SmeoIKQhdywe0BZS9dbbei9s7aBcTwWc5HbAkpYCGKHUC5ov5Qkp
/g/ssfaBDApBL9BzjFSSuh2kMmg4eXbTarYHg1Jvl+CroSuZm5jOv+cwblfKy9LRZN7yeSeHtEv/
Ye4kEZCLxrqQtXKmhRQoF5DhgNMCWaOyOJlMMAlqZo+yyEoxs+mMSjNTZfGl6eAz925/L74MhBqK
qIa4LYZrhkSzbsCRFXz2iIH6E8216cUe5ZSk3um+chwiHof45wilTEMyTczP9aay/RAUVjpsbcN7
/a9fvhL2AqA2/rUEvCkch4XLAN99LxZCgTDI3PnEEucrXrUkhoSs7unmRQsFn2N3NyAF9sjL88gm
lVVWMb9Rc9OUmUCNHOH7MT6Xz5wS9LrIOzVGgPTHW78nnDFbe4JiXG+7/Dzj3IsKqqXEoHJurSJQ
NwXtE4xJKSx7ZmWfpW3Tl13fhGDSvhCxoEmVhCdHFYLFs3tVIkNcxaVqGKjwOpYhmxhFOQnhve3u
+utslBN1wHXxqObgs/tYun2zae4EiRu/0w4xN4sjv9Juu5nSuUGO/JqDliFli7I2vLDZaSDcbRL8
PnyV5C+IllyU9F2M9aG8+oDPZy1D5/AL3X7LCtokSJXC1K4mZgAodfsKRNO8aSo0lzaIVLV7bUJh
Iadwt6E05Oj/qC7mbHqp3vk8kicMX1G8iybRDsmpWhxje+/0GL8ka7Blqm5GxCv0qQhbwJ0/SiEA
+bvto0lIYe/MONYa0I26Y+KOyh4ybuI58eZtiEnFx09wzRvaSf1bogjsT/nWOLR+zgaEpU8TXFkH
G4NKjDv5wY5Rjz2BoUQmSvLbRbf99L071b/uTrnLroZrSjsScOKZ33b7Q8pz/NUXNfzsKyEJxwhK
pDsRpLmwHTfPnV2hvtPmjroUOSn6Wd0NlI38IHR3+MdnGraRIc0fMCc8gFNnxOb4v0BhF6nf6kLr
pvt96qlDbBuKqH4zKv7obpiDYRC03CCuVK5Gjb2daiMFmAER4/QeBpMOyFXlOzJTgQnTJZP03QZb
EZMuneqLCxDZlOHK5d5hngcd7Bw7MIrfI7oI8oH8n9w/xjaBOSLvPYHUCl3wRNgd3jybNQAX0Rfm
FjfsDRByb5Dmbb/ojui76DrWlywD9ghGtT0UQk/LJ+j8Hu8S9uV03+y7CTM5DUMWt4B9OA3VtRfP
MCK0FaMZ4uuX1AQhXVRfB+J69Lz2lDGgDzrwbgtsLrFhiQ7R8k+QOONYgqUQ9sNinlKv3d/VepI4
nJj9mf3L/liMgZA6gxaPA81QJWbo+EA0PjmRLRh4dGbSv3DHsNNUMOdl/vVsyiZwEROInJmdnVq8
pPgbhj5bh7PNWZlMTax44IOYUxW/nXGgwXbwuSpNCLnaBqirVhkrP+ljbWhiwX3L+Egy5lcze/u5
nj5RxuSB0iK6NFeeE3jeakg+vCa3pZZI9MkgJIPpnOOhqp6EHdfosacnCeotxFZWqKNcRn6v/D0n
KEc4103F4oVgFtmf7b6/55+E49nyQc//lgtuBbW4i/9Wi8yAD38KSJFF73hSOUHqdWXm0QVv3jeT
fEY/guYIoFGOxFQag4XDw6UrPNeQwUNOAGY6c1aIdkHcD13X20YJT7QDF/ETyp2OshoIKLlJY9wD
A2XxNBCncsaK1Ylyp0RpU+B0f3Yg2WvbKAUq/AhRFm8kCQBxJXxuwfpK4tjwlEB6ZTJJxfypbPoV
wpYlP2BXEzg5Gwl+1Zlk6f3I5oKYbCQ3WEYdn38jz8lx7Ycrd+hVQZmpwXKCx7eRbibUjpkNi8k6
GsapaSY4+5MtECjFXaLKyHO05RFIQB1QvvkXle72ZORH8h/4K3a9RgFGo4u3PcSRSNNyop+cRI0T
OZwgXjljIu65+ftaQVIdN26YCzWQP0LG22XEBAg1Yptj0zJKer3jMX/xLY4n5bVu2gsjbYLShVN/
llwTsbXkTcqVUzK+6AiV/mGKVEfm/AYJXb3QGcPs1dpLRcqM+LOiVe0LC7SmH7T59ncah0N2Ib64
p+QusbXSQz3CrMJuNfab+jY52RS3oSPZVWea0lE9BRmdGIyt9xFmovHubtNumJ5Fm8dcXAcsqFBu
ArVIkDmdfO57GbEKIVc9nL5Q6/rF15xTXSswUDY2lk8I3hmBl1kJZ6T1AoHUZUNW/tD+53QSeTR1
oV/nfEBiHTx17yChzKslRZ3/3UPG5P3nXP12Siw9LYSwytZa46J8mchFkGzd73j9O6MmJhwE+Qi5
jHJAUVAAdzxgYmrW8ib6nR0GI5CeZORnStLODlkDplSrGOV176teI1sMafY41clxmfPcLP+8IEAa
np/KQ8Jh63rP+6itumDREmae+TBmjgt6J8xi8mdgFJUgu2N47cFTZvrR6Pw78sCXfdtICIgaqFnJ
OXPR/DegbH6lYUPhNiiXvEbEE1GmMyUkzSjWAESNQ2fjJtNiYPPWFMJNBBbIHtCqR/BFeMKvpEFR
eXbd0EXzoB0zLPRG79sbk3Yc6yo6L6+pBi2z4qi2Az5MmXKiMz0NntOx3AoIwc8tI6GmHPvmywqK
2tJvP25XjdJvOIs39zVkcDaPJ0RLtst+soU94BudGdv3NhK0MeLk7WSBEXdzI9JvcTMN1U3TGe3a
R35sKoGydCe+mgyfaLyNEm5wsXOFWLSOXdrvHogYFU8pr/ZUJIjZIqOTuX5/yiyOHC2XsesfZjbs
O041KNt3ZocSk327f7MGXp6jKhYbe+a+VIe/UMnKnzc9Tq/KuoE3jQ9jr6CVDhiyZa+ZqsPQzu3c
HUj2gPA0f92Gu+7mizAK7fEBVnKRabQnckC1zkO1/mc/GLgmzf6Ie+gcK+YOrMvPpG9j/BGTE/j7
CZJCjAKXycL5KMRTTv3aX8b23++vIleWqiGueAHg32o3gv5E2q8GuqZRpE+apSCbXcwMSOUyl2u3
VWsGyuwS7U3FQ8p4htVjfvSMZf3kZosRizViJTummfuki+uRLcK/IvLihOHPhTWiXEhMKg1yeg5R
w0zMmuud6E50wkMTtXVjdWmyihTS+qG0rpOl336daEehKavOfLN3dsJA3m3usR30j7dP5jrp7KJ9
2AQ+CKILgrkRY0WuJwdc+HMJE+yTB9VWb1As3WNTmpZTxEnusdH1ubJvzbateuqhxg5r8Rh/6OOY
zvBUin/gxKNYOhHIsPyVndv24issBr1N93iA1kdx/EzzGZSe7hCu9WKcZf2AhwZXoqzvz3/cGCau
zvrLtR0tr7NaMznkQFcajC6P91792vdEGm35yt0PSxSK7P0F8x2a7BvJp4d3db108rFYuh1OtAex
VtEDjFDV+c4ANoSWOsIzHR+UQu4O4nY2trsUalikSX5H3LOyoDw3wBwqsw1JF2Gulhzr70iVAp4E
/LGi1G1hZVKIuZUg7MBvww68lgsGTaolo8cy0aE6YJN3zMbOrNWdI0lvrez8jXBTwU8rmLrJVUrR
ObK06zUk4fDFuQyZdoMTbJrwDB7zBliCIaN7g5RlN50jd8QLmnmAsUo43gM9SYE0ZZV3jFi1CKMy
xf8b3HHOBRh7TyICuozJx5rofSBA74gX2/VidVKXNw84xDaXB9gSfTWRR1E62U0k1cmUAirrQWlg
ssg4QUDVitf1MHRdi3owYW9TKlc9fxhYpx8z3RV5Y4+rqjoZkfMnU7pmgGiosM+G8Qbq7eRaBxQQ
0bKgc8J675+IjxnNlGh3b3W3KmoYWDUS4fRScbt9sFRyD3ZTL/7N26lIylLLh1HqECmJTL4qWRAZ
xXz17xI3Adhtqq6L0msW+jZTOyK88DGye6cPFywKGe9lW+MKGDyCH4LtwV9TidAZGiwDHvjByXiu
SisJRKf7tjxmZuV225o11Fta1FxO0618MzlvAW5IRZSYwy1+nwHuk7aLvh7jVoFJnJu+H5RW5NzJ
6juZFKJrwnDwd+Zc0NvgScqov0XDgpa0HIyVF7C21dPzOA1+rGDZsQ0IB7iA4UtPBJrbCSr2p9Ei
v29HrTQp5nsJhYd1PQIpqNk3S+4uGXwokCWKSf8OgbxrPQvcEl2L0Y2Cp3DTkww8DmHz0WSf8XDd
xzldc2gHXPV/M2hv1ZZrLQ7bWKP0F8hRj73g2a6sTARk8YfwHgBYSoQ1WwzyHHM4i2R9CRhK+Cxm
gSFhoyod1CfieFkSB4M1sd+icJQexzGzZvfdElS0Fe6AaNhws+yzk6+8/zS9uZemiK2MXIaw1zYV
mbGxohq54cVJz+xMkhJTe1VKKnOzJslaBak6FZ37h7jWcGhyX/IhAGs+13b9nYsaz5oX40gccP0M
UZPvbmA7Zp65wKfhn6gmi+S5A9xrRttxQ6X7lc2s1BLkc0od0tDhCv4USv+VjLaOcxUIL5iyzEgS
4qsTQs4YUBgRAODvHZZO/dAhGwWvB4Fhc+daflhoVppgQ3RZwQ+CnDq1kl+pynrxmoWM7aFcE+ay
D7XopWDNclhl3BUKOKXEsKPcUvuZ5skF5F6lHpwFMKDQjxJRd+yzteRPkNduslv3ANV11doX+Qkc
1f9xCCSrdjPWZbTPbI8mNF//drSl5idgoue6eXDTI5i6e9Fy9bDRWjxSVxnoSQni8hY961l1+Su0
rb/2UNdLE5QxXkZdyCNBNH/juPLTQCjz1bF1DhteTfRZigBEXhRKG4ccd2fNU6y+HjU81sVtQJ0p
xxq+lPUJg8oE7wUpKv5lFNuuM4MVh8iv8Bi/f1AmsY8HTBeFf4KuAZT7JpKIhSOSc5/+jlKF4nHc
7rwS6pX8muQxmxP1jaxVin1i+jd8Wr2eV/NiIOlxv07FiceNefDDRxhwQY034RThaiXfHBreFN+7
SywP7wxk6uzwrungr8BmpMKypQgvDQ3FDecdfPB5xCsxtrPEVsiqSfb9wphYH+LihgAk0xY0yBJs
KdNddtKd9d8hc2m1VwNSRDvIaRtwDqgZVv2mF6gbWW0qY0WG5T6GaxwOMlGOHoL2yZ5gRsrQDQwx
hDVUdDbtMYeuhO4PYSkS73T6fnWNux4muzuruiOAR7vef9riCmy7gzkUbDgblCfqkzmGx1PKWrem
wL6UayieNJKY3qftYXTGz4cjNObRHFSjep4eKwiqPxCff76IsKQ3tVBhx+psrvINtemv3oOwucY8
lGwapbnglWfiofiE6j+PABuTVZUZHk0R79yvXQqRmbwworodMR7ELJ6nqsSZgftgsqU3A0ows/1k
zwdhPbdqoBMbYZKMWpl/Hgt6BpaUREEo0aTut7iiLAmkj4QTHip9MKXDOB66pd48QQ9Zai7sEDG/
cHSUKFQ6Jelk8vIyuC2iwvdj83J+TsUj+UPLv8KNRkqujwxy1F1GQe+Ak2xsLLQT1QXjVFU4SZp8
Z/NtO1HKNROviXBnEFN6QS5rE9mEQ6biHXtAvyBkP4K4DSbLp4xcaQbQiyJOZKwhz6KBqaiVA1GE
/tOMJ8kEPnH7XEEMTr85dQMn9VFKK14fdEOeZ0z9GiQVcLDA2jXTzysrxIK4VacTmRTHVegcALOn
5Eodg/T2BWCrECR0LIc9RySfvCh6YGDoedGw1ZSmnkfF3caPrnEOW0lf9yPQbZUKhJFcg+K0j2Ce
htYUXAdq7qgJj2IImVs+c3RAsuRuJUaaN7EOcfcWv/CVnu50nSLqXwl/5v390JFIB5W5LVQSiKvY
OWhypxyyVRJr+QipPshiKCHdGcYIu0Bjpa8GGupHLHUnL6JpeXMO2woQ8PN0fNVxKVIzsLHlIzAz
TK7riKTjoUR0vxXUXwghvapyJ4MJIoW0z/E1daDJ62pV4xw6yQe0rsfTkwwq/hYq4SXrA9qTBbzn
xyjyIl9DYmD3T79EUFUkw6ojpY36RmoWi2BT6A6jSXLXBlWGciLD6M4AMhkiiy8Qa+54m+o1VMqg
grHPfgzevFm0ycYk6+Gr/ZEHgOYXWm+alA0dk/GR24FX44YkhokwwUQ7AeLyFEP4BZ5bidbNqWS9
RgkOBRnRprU/6vkJi1Vdu6XykOfrQQ3mv5gNazKFsaBijfe7yTU+74nBESXQvTDsoeDqAVIPeGN+
yUN+IGEjWeGWfF0WE8ox5e63wjlX/OZR+bW4A5KUgYT7+n/Rhr7saegGJOvKxdR1KzRpxmccfA6Z
fVOgRSyMuyrroLHIc78ET5Ghl83+AoZJPMJYWJfRluVFMxakghxhpY0sCMz8fkS01R+7uWftVCJE
E467cWC3Xt44zmrTg/InXWVp0Qj6od9BAlZSDmN6Z+RPTA44PyNZKkpxlSbz6JUZnsENPHkOourr
SWMALvapae4KPobOQkex1MT68I46h8yB1tT4TEAQYkNYHEu4TqpwkZd1CRh5BKa52cEitzaRthbl
C7mU7QErShoDHRYzdiyKkrrT+zOSnLa0HTxAc2Rg2SkTDafjXzkBl76fCcXTrQ9M0WuHs3CaekhD
rho5Fnw3QjsuQWsrk6C8sKsJ732WmNfK35zuN0ZuInXZADwRzSQ+Rw6py73Io+x0d/xpsK2k5jHH
pu0iLXDUYpgoSz6tnmLO0OEmbIOAJma9R71Zz4hGHrOGA8hI8yeD34F/QcWdSF2bZp/uQTZatAfh
OzCRpV0cykNkO64W2qcoOQg2yHPe7x+tmOVsw+OS4/WWyCV9e3hOh/2ZCNImsJagUETgSKy/ksC0
S1r7t8n1fMCG8U0aYJtrbKJbdCe+ukeja7+vlGrasjl/8vey90yUGtSgLQtl3YUOrK0SpKvM9/+0
07cQG5owuBvsyVewc5yypnMf3fo3L9e6NwopfAaqLafdcqUSKQTbdC5pSnyIQwtd7LcbQjgTJi5w
SLCFwcO1SEbuEA8gT/JnUo0XYxXWSOvRG5KRIKf4Ysdj7WodxSGyiLwcbYorHJHzwjz+JT82GOOj
k1Nx8+BaAaEx0sKoDwsUB3OsZxLoLLmL5ZcMpMkXrwZpOSq0eizeqPyZ62PVk9hvb0YzXA7fnJiQ
xynDOQI8cuRxuhO6L3Pg+UqdCbQqrVOUubZwyGa6MCnMx3beEt2LItZZQ85CMX/h8TZL21YZXZSw
u0xzDqyGQgx6KzRtvgWjRUZn9VVZ654ieXqLLr7kDX7AeE7F+GnC4PlZjf9dA12rev51lwNm4O13
8y0J3r42PUYPV7vfLMCJNUc0DhXOoB1jf3MoxtiNfWhKmoC+/Q/J92Y3A6MG8lV0W805K6ZwCxNo
9i4BaVD0OKrZ00wOA89qzx1clFyX68LaQvU4e2d9aE/NMUT8j4GmNRgQRaJeJ3YDgPVL37BDsz+z
9T2S7rzNAPTzM/7uYl7dJ4DZ1c+iPGfOcPheXhQ+ezI7QJKC/QMJYwK9zcvYXm/IPxxUDY7tLJS8
VwOvpA/+6+ziv59UoCgUUGcHcdRkOR4mGnyPjv7lYmRtdrdTeiHYAuBTVEX9smbFQ4y22x6LWynI
aPyGe3G20x0Kelo2geo9z6UBsr5SoqFbAN+JbM8BjCd3c0nFouGlUhSgvtyTSMP4jsKQHhBm9lD0
/8RgDgjBUfgr/LK4iuENolqihEY5pr5a+xNHC8YG1DI+ucBWH3GfmsIfpFRyI2cYzNQ/rVBt0qxB
DPFu9s5qq2maidaq+NTC5qIA/AZ2pv0fb0UpIRWj8JcH144HWdfH3NKDjnvfqylJq0FyxViRABHD
eZi700gTdF/csVWleTnuK4CgI9//KjAXWfjyk40RCUdJsCuica6hnSOea0BJOoV+RizClG2gxnXa
RWM/XSGxasMX5GsWshEO1OXbswjqycTxv4Z4gK1evfu6tR5M4272XitD2AZaF/doayPMoahkp5Df
VIQuXxhfBYshJVeWA5Z70g3/83Eal9ISk6AxoQnJU4rFe0gapIIxzfu0zMLgTDnu+FGxRaTmEMWe
u0rnxODj9u9mqUomRxFJ1H4RuSQ85KvQ0ndJMKvFLE1hQ4zuCb5bneSr+pYJO8bgk+dZM9utH4nQ
nm+uZ37MAycdDvGLzK/FyPAVQmsNIvlFyWhFlW80ieBIkwyMh+Kdvl24LHc8oVSetjjiDkBVLoR5
29dModT8vbDWPvsvb3burxBkop10ZeKi7QGytSH7UVf75PaGTvMZWzOJDYJF2EpFi8E54HlqMhx8
HJ8fNwPltXnncaaowugfgvYH4z6gYevBHxPwnzjrDvcuF0Z+YUez6l6TLuQyA7Pl7RETwWF34I9b
AJZaAIKO34vzXWmkQ4/dlD2OF1G1o/EjPgdOGg78zR5FbNqXkHBUKxLa27Do2sgIPAVHYLDPy3dq
q8CSEnotoQMTR1JnHRT5TWIds62L/3Vcz/PeukUSZ7V4+hODim5aLH+sfoUu6zgYL877LQnIK3sb
MugnBadC0MjoawexwqvMDGM6uzrZdszdBNeI9TZKGwjqOiGLvFE7nXuvCbE27lKb2u26E1tYWye1
g+ZJCbZ5O88bOCjbs3aKREXor7X1xv33Squm3Ozn5xWiabQwznws4L+MFgNwZWxmwGrQqo5t+ih7
v4bHUG+XQqzq9QIk2kKGtegouhIyio/0FPWwkWYy9JT8LGPDzldquFibgnODxod2Y9xjEW7/QZjQ
1DiemqPtLo5uZFlKjHUSDP5aa1B5lK0R4B95v0yT2dd3o2p6Ul0vAi2ccD4OfCnC/as8d0w9XeuG
v/0lwZaDMsapz0dsl0ZH/eFcwHJ6uMBBWeLj2/p8/1eL8ArQSEyP9AOszIUhFZPKZK1YeUUY0Nu9
kU4ktiRM6HJjjzPkesuvAC/He2g5pyApRdTGVgtvqlJ9b2KCkmeQ2Y1Mj/t666yyRAe+VHlnWji6
eXzwxJ8nxiRRdEOmb6/Ut+drFoyWx1OFwdZFOXHvTYJEu4IapbdPRsXdc8EtGMrckdEsGl8b5UQ2
fGfM+v9+BtritRtJHOTONycr6yI1DXBXaxFTTMTJvIkAwJqEMm9Vr+8M1IKIoRHWRPHPLvJHPtVk
Jwt4zWky0i+meGz87VRXMM7vV/0RGUfOg5oQtJMnU84cN8KDeykIld1g9eE7NyTqGilM2+1eqZHo
VRcgAVmVQBMCyyE+++POPlw7CaErFvTXRFmhIXXr+5fpnu6sUfB8SkfE0uDhazbBevXktEQaXjzn
URRe5h+diw7gLjW7K7epwXTLR+ahJMeUCCxzBfABTVUMXhMkGMjHprBjQ4SGLIavcESVv7KJKcg5
y2fbubBTxjOS9UNV/2S124GOOYy3jD7Ws33wDRUN/QRPY3V79nVAxcsG2QU5L7cDq0J5qPs3PVKm
jKGfV1iUGTyzvSWyYdXMVAe6l6ixFhC1I9TEh/ISbq6xD9c2B8RGz0cufWoAZ0xAtLOrrWgd6GPZ
dKd9uCIauYXR7P/pPW17/FcJx7zN9/4wcolJUfbsliufO38TdhV8Hor6scLcdKZfPelzj5nT9klz
Zl05yH7xLj65ePhIvnujFQCztvSYISJN4VnIMFA5r3rJ7IOwyAE4guZBmBFp0nSMuZ+JFesPXfmG
rZFlJVatbZ4vh2IFGJL6wfc0bRm6xWeSk07nxqk2hbw9vmQiZyB9n7tDagL6EwuNrf2FDgEsB6fi
kju+mkZIzaP4zhmv4PZV0brNKwCui3UWilAGManODGtcDEwmdd6ShVbDMlyPqxivnqovpw1q00l2
2m8SzXZ8ZFzdVS3zHUy6RS8Uj/HeTWGJTQUMLRCMsWY0VBpWsXh20hffnvCSDHpIaWaPSneRND3e
LuncgqsL0cPGgo60OqliemKn0gB8LI4k8bBVt7dVeo7ssbFd9DP8Ojzdke7e97LZpdn0ExjhI2NQ
WXgVPX2fmcUfZzjs3YcHJd+5NfOIX+8GAGJ1zjQZpSu8i3ATFFU890vFPRQzG7eLXt4T/3nFGaSV
XUXx/jXQgSpT/iximq4QjzmatWPR9xsBldrM7PnafDNYYc/Dqru+mnbNT+oyb8cgs18vzKm24xZ7
//qcKv767yisRs+Hka+Xg1e8zxwqwPZ39IH34f/pI9lC4Lk/7A1xvTQsQWfxIaIwQdeQDOli/sk2
zqei/Wd3tLA02Kw088wf3c34SBSzHTT3BJtkq6nEJPVxuWUt+kX2NcJ0WPQOWdpc70tlqRwRkpWC
ddGAdtzrCdW0zKn9tuEJsTRd9FHtpzAsUkR/9pDjRu6vmadKBrle5MhNL2Oy6E0RxEjw+YmVIo8N
k/JnKD2JuCcczalO/G563s4E5ppoDZh9kISA1oLhgs5S412Fl4e0fIVg+A+ytt9HcZCxLKinZ+EZ
YdmEqzIk9L1gfxluHrvxByytHxK2/bmHfCWoOr963z0ehYLtTVTmRGikKfTcLDyilpWd5PGbyhGT
F6lnHt7lqLUPLEqJRh/+++WiW2RFNRm3ZjFWVcvVbxQwOvXx+HHUVFipsfcZlKtPueM+MRLsRtnG
hA48glbRgeHAz5oeA8r2ExYhUKt553YoGW75p90cu9zFXSYuq8E3rRt9MrWF9nDNSqu05H0ztjhF
5fhOMPp9YMNZGSkz5hWbs8EptEG9pfpXbCK7PDGqVEf2XKValuL3tmUhlN0KkLBo/sqGzpe++H8Z
dm1csKRz40xRGwwZ+wng+Rmm65Hmd135q9yXYdy8rCR+iwz3wT31lRzKdyURU2edg//aPklF9jU1
ElbR7Q/9m87uT3IVuILjiZs6ztfZD+3TvmPDBC0tU29Vm1UcVvv3hyAUJPDQJfLGLi6g+WAGZBcb
1rrEbNa+L9ctKaByUBMy6BQpUulrwb36/Nylai5zP2thvX3CPFMXh6zeD82ligbR+UD4fCVvmxuY
7kAupJlOClrvpGywf/H8eKsAOW+uqO/LJkGiTP+ToS3tLhHy/J8DrS/k2c+vDCcyu9E9oKETuMLx
D+pcQZZP/pXuMCD8tuEbP2UuaA8haHmwBD+La1c0EsDLzJUvxKBkboRQW05pn5nOluXwMu1F7gEq
3j5grBkaYepEfoHpRFZyHhAxfGCt6mhhoHdLrlzCnwW/RLr1k3BYRKA+5rYWDFRWKpcU3Fz9BCjz
jf9HirYdWWrANTSmH6DLP3ESSr1qDMtcoHcUKw8u0DHX8R+f868T4g6Evi5ItK6uQ8B8oZE3hAby
ac+JamlPPzMRDjpe923qmDfuBlZ83kgeylwliSDSzY6tx6GH5E2aMG5/mFX5f6+XMkFdoCaUsj6J
Lqlzf8pFBwpmVjB/iHGI2ALqDdxBaSNmiddDAYpT2ZBnwLzPZfCP4pp+WieP4YhCJzB4piuKVlNy
aYPJshQ4D14Y20b+LmuPf1K1FwY1bZ0s0Zkx5egrHBZgDEGSm9T8XVZy2xMmiA9+T2vZqqLl4lKg
Qqm+W3jOicueUnP7HQNDXnXl05GYMK5dPhEoXII59dp4FrlPE3a1D3OWc+ApTpXpTkZN6ZpJmeIk
z5HW6PzBJAIOTv/0lgdrop6v/8k+0lmv29m6UP1uc3elGBlTeQrvlHMUgbGb2Ly/yqfWAWBUZtk0
xdsviMSEdarsyIcJblBrl2GqrpGd0nLQECqAoN6dcFjDt8Q+fJqjAcohVc4N0lfB8DmtPnlfizJ+
HB3im2LMUs6H4UxkGupVr7RwHMYIBBNzDYdH6Ce41CtBHVUkbeJReAPAffGlm4u4GpdZ+YXR+01Q
+iCzg5HjGFSzpf2bWS0X5PDJRnSbWJGhXakNqlpynZ3Z12NpieBPHrQeS3DSceZ9mXwN/jzX+NHH
KPRUZjOhBwq1Hmw6QaNu3FbOrtXrT7P+9Yw3lnp9x6e7//IrxoVRI8HEFjTpjuousoIOtOimtBxz
hfbRldDc7uhpN41WOFvfcyCIzoUHz0Fn35zkIUfQRreDI+ToWhMDYurdE+mffg0wVXeQDLjtny3A
nnMFGaP3z6Hk7cYaRhsXBt1ZSmI9+m7cgeJadrtstnReSfr0qtcOMa+UwVTDUvSy/LxMAATteatI
sgpkYkALGI75xIPI0IsqvT+m/XSfb8R9fcJdSSOE3TEmYSlsLDKrzt4Hp5Cu05RXh0c0o1Kksu/0
yROUgwEy08UmNo0Bi9dcN+e195GieBaUrRjIE/M93kQ9DM2bp7MtsjNwFiVGusLW+Y/eTTImYNlZ
i5foOpq22CY0ojGwaHJzhQv/SjlDfBG7B2qLacRd5hVbVVKLnDlLQ4iZB9dEz0WHgnT5LWnfqyPv
8jvsV/NYOkx0QDv9Z2LYtsCfJbqmoC7jY7vOquBqqGvHb1j7dTyHhv3AhwWqsi3aNxfu/y2Je3Hn
RWx2emplr/V5ZSi5yVryZjd+olzbt9rXB4zyk8ZH5NjnRpCtF06vmk9RV52VPB30tTA2SyH3M0f8
zOVkUcwo+gyQ6BLZtn2n/8x9dA65a8v8pjF3+1MONf+tqNEy73ItlY6X2vDOzAWamI6m1Qsx+4gI
i+qoTTytn6JRRMD0IDiF/czFN8g4jnMqbcsrGmAalUi6p97FDMCtXlHDXqewZLOYG6i7AvEwews+
x3OTfSs/JN2HOJj8uZUvoefHnphPlgJGFs3biDuh6N5zWY6ksei/nXTvz3h0SoEdsQhFm8kN+pGC
tzrG/HVnbEu3J18KImpGeEWsyLTiWGdwyDFyQukDjb2Y0CXg3w59no/VM2QvXdq453a7qLIGdmN2
Cc+ESKW1D8MGVKu2IsbfeaJKbIFt+36tqxGxXj4wAEBjUgeX7DCDNXiWfcOoLD29IBeHNoLVcmFJ
lAjTmd1LeYT4UHyIhsQrllhrZNPNMCKswMpz+i1Nik0sSXnEqg6EsPjn6vSR1h71anF6sr1W8eAw
FhnSBKDTVCcZdeBCsTCYA/vuTudnu5d9ZTmMiCXNpFqFcHj4I6aXcWQ2KgxRRn7x28nNsE9FLrQ6
LNxbb2mJcNt9USbbR50tUyrdcbqAmaETxhCxj+Nk6cCmTR/sDzmygBOuvEqNxxfOVR1PAalI60c1
IDRbCGesAGCMdS+5L4wZJfZ/V65mWQtE6EqeigQk+M0l7nyA7zVGduowT/okhXVVa1BXCQo1b6tZ
v0r6fo71+V+VuU56bbe+AU36+W1WSk6uKedX+xhw1yyivoMKoWNhnLQRu36Ahf+eCW7xcnjaS3Uv
nJZoQsdsa7ZJ4oqCHRP9sfz8eY6ZJBV03+brZFLu+ZERfMxrafXMhCyEG/JsAxTNVYMwkUSLCiJ2
4t+AISEEuTmLKSMFHPHMNNl9du18qwikSVExUWCzV5TCDekyozm/joNx8/4GS99ngOBIIQqDQliq
iUTMf3iXJW7fQ+j/WZERwH0MitPEcXjAdQk0w7QQxDsJvueVnKcJQm4VZ+hHA/kW/ohVCEsne7xc
befdcCdP9ltJGYWzFmgUfJAMvsR61gnmFdwWEacA3k8XXQpaXFfr84VqTpxn/Vxlh5aw6UVG2pV0
ibzaxs2CCZOBi3vnF2jLvw4W/A3yoF+UUqsxAYsNHZQd1aWRwCbGkqinbpAT5brSpfRA4Fachd4T
kBxfz4GwOnAnNy+tmtfrREtHRrjP7i6HzRMBRxXATadBnnjsOMxMg78cK1jUQdAl2uCfI8wGCyXS
vPKhWYUKypoUtS66/rTSBsMf0C74tlYmMZqmeZcgO+UVYPNJBw6GMsEqLi6mtfIwrvcubkhzD2bt
nd4mpv+SjsQMwebJZlNHN8XsXHvLYcUCpt/7fnfnlx+y2fqBphN73i7pbf3aX5vd5aISkTIkzBU2
nTCS1CeEZ9SJz2JBHi8IazHDkZJswq/HrOph677OISLUXs1K3F1vw9Y7Tx14Qpimn/xdJkcqGxMs
xkTtTd+gxe1IpX7EsTBhRMDJolOa1ShDsucuvAzwdkz5vVtMDrpprPr86hlgyLIH0fcbsNEQIS2F
1QiKJbapxDkkEA+qJGPDknPTVtXj/ywPdJVfa2Jgnhmg3DVYTFOZg/XxZHsyZTP7jzGkMe7N5Wms
b7PoBjz4EnOq+IkyTnxi1K2m/PH06bSLlzpIJ/JcsIwIrqhhE88N1NK9WvdZqx47lLcKeza4padS
XJWN8mzsA6KKFgzGbqZNfcdHIvP7AShTIlvwVk6x+3rs8TD8AokcmFSqEPHbLX4mhtbNoqAZSAFc
6F2vGAoQOjE7jF6ZRrL6bCCCCztC5K3ZiLNG7emDqt4v/OTOiDftLEUy+I5WFNTmPO/i0Tyjo3u6
WcgVRXVvBENQkYgt5ToUtRNiuWG8dZvs464k11/at3ALU/PiviVALTJb2DeLKD+CNDetoWlvgC4W
HQJAP9nNcrq6vCsy8hDIASCu+CbVilNuQx4v12hyIPdrq/WD8VZ7Coruc+TmspiFSfvDAY22MNiI
JRFZiS7YXEcdrZJ4AyASAD6ZONeHppSeSwHJ25JDqDhWIvWwrmZ/p14lSACp0W54xT1Pq3Synqfx
w4E/pEkaZmunRfu4+HK9yYGsNWGT4DCbYcHoKQPx0xfj8egDj/6c5Hk31z2zZUzuqB4aFfYY4Wiu
m48/OTXW8olv1G+UoFWeIQZj8/nQwERqPalJqdNe/nQXQ0aXxwTztbVlVfK2mtOb8etnGW9YyvTE
i2al03lKaMAOHmExtx1cMWs/DfDIqB1fNalQzI9LJPe3mQlMrbs83JGQF8vuFQXt6uY/1rO5nR5V
kH5d36TwJh1dt9hEv7n6ihsE2Z5+TXDaJ72ch/BODhGYRtsFA6sm+ZdTSodvkficj6LO0XW0plDl
h1SePQtrnoBE4DjAYSziC0Ayt6E2BHuz5zC38xetAS6YNlhZrGdF5CqoRwe+r1eioNTiQcbTvo0Y
0PGzwXzo8jf1gkxf4VaO79C8Se3/cX6qypgyehcGQcM8/U+PfWAbKcSXQuIOjetX3hN78bzOwAkR
NQk/XQ3JLGSutugWhsmQN03BsaL1M+/+e32h8VYv8y2KZoTPAd2Khc2KkhbtWZlvCkzMhBvRFhOs
lQIwGqChmdd+WsMuoua+XSjAJKRvsBSacQIdDwshTgE2sC8uodc/u0g78mYy7bN5gVDeEJ3BSaQj
USzp0JalNPpEqCf22kThu2vIIJjm0t977ZBvbuxQf42LoltMFDkYpXNarKUOAj9qQc5zKFBe6ctu
a/HltZtQeD1kgdBUAoiD4qpwJQFVmjUvx+Va58hOSEJ2bvWsX3w9o3Jzi601YSQHIWq0rk9LRb/S
4oJ8HnF6yLRVexioSb1kDXz4G1ajnpY5gFH2MZkHcK3oiCzAOgjfgZTYkPy5VS4XLOW4bEmFkUT3
mRLNuMKv/RyEMILkl/RaMW0zNrDzz0wyn8vslg5Mg2dD2unvwxiJhatUlmBqLEqXa9ODlpZaT9Xx
Xj3EvRPQfqdoqswAak1sAxQw2DPsRMpee2Gv6bp0dqCV2zmXvFpy/1rLmkD4XOJZEjp8k7B3fFD5
qo4ZMOapwHxkATyaQb7tXyIGP9MY/WiGkvs7ERP8SyfwPjcc3rS0A9NWOonLcYJ9/yRRDR7xwknc
3JlgOmVcV7zYBmdr7G1AFVRp3PRQE1FhFbTdVFvArnrTqVfFZPaBlUvxQFZkurwgEV/9bcmVqTFa
qd9uw3TdFXhtmWXqpnyhe3DMPxwynb6nQkaP94+dL6umAWeNTngullVye2TsOTUKuf3lFHcDXanv
09PILub2YbA17LVLYCsvJbAhbC85nCeeh98UfcN/i5fQiEB6MorhjX6ueKVyaQxZF1nlnFpmovoj
ukBI4LAPCo+S/xxLK/HGm7m2Zrt5ca3pEwQADLBBgPzIAkULEVbtcxOXKSQXgNbUKYN3Be7xCd/6
nRpWPjRNIcUFmzghHHJbn66zulv9WcIV9wpfm4fpxOUkTkbsGuzDGPP62Ut8oz9O6JRo0bCsokEb
dpEKT1SAKZtmSM+Zp9hZaW7bzlXyDXIqma6vNHAyXryGe+RM9RjjCN4HGCANI+T+nI1peJl6RFo1
4xd4yFfK5sjDF9Ep+fs6r8+y6GDIoN+oLWxgp6Xz5R9qBuIqTiG3s9rCfxUEwcsGQQOLw7UNetdW
7hwcN4/opUqZWWnNDaliBjVOYSfcW3jRRTkLdWDx1amf+XR8aBNnr8fze/UuaszCUHCOb3Cnf00U
y4sIiVu7SKwcVIWuOjlFLJ+WwrRVSchauffxRbChHsBC4+F0RwuTif7hNYoZlVDGiwI/uJ3lzpPm
7uUtKp5/RjsoX6EudECvOi6tpX0dEg5yE9f78PWBeYNMiIhIEylqVQNyVdKDSmD3PzQgmL0eqp1J
FrdletQdJ5rn0o4wcAkIkS1HykrNKybNbdPm2MOXCQexk6PYej9M91LHeQFzYaTexTU5OYEzCSQi
E2Idk4drlGOunVvbNN1EorrYz+sRvJ8vKv4sTHJErw17aYkAajAnV+VOHhjA7v2bI/pFUKG6rjKf
AJI0J+K777mmw6yL+uMNeweDWRLPf72VTqDE0iV6ESp4p5CfR96S+8db50pegd/wRl2a+eqNrL0W
U3cYoA10uQFivdiJLQmArhy2+f3nJN0U5g/YdASPwZq00dxgXmq8AkrYRrN+DFbQqdqxy9hjo2mP
iMFJ0hIkgHT+sVuBDxuLYADXM7F43n4/XKIjsvK/F+OkDgR6c0gGvsRGZ319OJwrTD++G/aqlSi9
amU1QLXT76sUifwsVql75Tp4ih0LrD6sNm5vp0XR2iEMQrp6ZDv1txoMqnKYudknQMFx9iOHi60F
u5ZDkx0jevuEIw8EuCDzCbFJ+u2s/eMW4pDPKuGzmny/I5qzVo63DB3lQsthRePpqh4gMPcPscMI
dw07uZBCc1aHuwKpQmaMV2+zTrB/h4ASXfL5L5GtqmOJkeomvnju5ewInj5YcYvsxl+0AekTziI9
XyfjBnNdnuLG1HQNIG3Sr2YL/UqQ27b992WwUD4TEo+v5uX6j+q2Wtfa/nwWAgzkH1Qp12+Ew9DG
9BNZyr00WEokT5cOHQlJQWuYxiv9o6s5wCl5b6hVLfwSvS/PLvl9ZeUtPvB4YqyY2Bm83UeIwLOQ
MXqwnbPbDI29Av7JfrwwkmzZu2NvFVpKk6IS6yQ7+QhGIegpT30uJAu9ZVNi7mUlO5z3ascuirME
rbkaItDPmCPitpfa6jnkxRMY69XB7awkU/CBJmT/ehDh5A0enwmiDCjYdtBydScXr85NsksC8wZ9
Ysa4seC+C7Ellz8timsV+2yZ5k8Kc+YGbqO5+5yqWYw0PCzAMR5CCFEZSiHdgCWSfI4JMhX15MYf
FmG2C1w1riBmA1DukyNnpZW/2ACZlUOZ5/xpyGVdjkhxt8pOY2OGcV8e2CvJyjIhp0ReH124m8gK
d32n7cdfrqNkJdCIaGGgNXcG1+WO+Kn1WOgcRevIV8BKCJR/qyD8AAI9b8PyvseXDrl137nDrtFZ
BlxC0NBasst5SQPebxze0so/+2h3REt6IO6SnXQapnXYSxEjUgwHuJnBZ3Ej5wGeotl2ekETWBGI
VbDUBu7jRZ7+yXglB9GgHS7a9bA93u+Xza7r+okfnxpObvlAz1NEV5sW5pWY41L+MYLM9+ZyMk0O
5TAmW7+BKHJ4qcS/4DLGdB3oZ5JsoUul6+WtPJ8tlp3ffp/N61bi/Un+YC74sUcK1uyzs9w0ihpA
FtuX9UrrmdLDmi4In0PgMtZS2WDnjeQU3CI4QDLTnDa1XLDMIHUgJNf3RMoA32up9Uo1C8ZQ3Cl6
7ywdznvbk5As58q8qRjsIMPzFehKUTeXB3+qXWfFLbBPSAIjhzM5CZCPbUcEnexJGJNuM3hU6ahA
7KZFEBfsWucpg8lf0SXVw2xgjfWdJfrWiedhYPP4T/Iu5UlfwZxLrWqW14JrxmCf2pPTN9IP5Hxt
euxCSS0vpZhY+oooBK9z6GT8js5/kNse1qMVxxE6txANaMcx8jJw6N5NeKzsxbO6n9K6PoxAB4Qu
Irhd0ON0IP3yFHAXthe208Hr9BnYC04Vze3EGMzAxXEkbEWT41MIK9ibhdL/UFtJw/vcVeUm/EwW
2DGljzlPShmmau5VHgVQIcXzbtpJsSbNYybv6Dkxuf2jtlqxSZVCQqXKPLem+MnI+eyx9iHZ5i/f
UtnyySrpZZ7xSo46RNrfW8ykZrurD/SYMyULtwgc0vMms/h5Iv/UHBEiDg+ilV15GvCPo2EAvWKh
ZstokA5oE+GA6/r7xSGutIM8fiP5GtmtI27jKj5fgb4fdMDQOyAIH4qZedh6ZF65xgjAIIrAbhuq
RhgerWfCfbgUaPvn7xwqG9BibfZi7RfBYCgimknLQpRSc/3lyVatAyQ2FFbNXzFRhPChpKhGFGxy
T90V2NST7wTVQFEKALumQ0oBgTQohae+R0HFUfVNknWRLY4yxhcAKUmbHm9r1cMSTybsWGNbsiAi
1QGDHhK/p1edf55Q+/a/euYzzuD/YapkupkhuKAQdufQtTSvt++l7YdJcCfDfp0ma7aQCdmfsQnB
A8RDHa6K5/swye5NX7gZ4YMgFipgPPy49j4zW49xB7em9G3RUD7RDN1rlARE7Rrd7xtr+u4NClXA
t/1SSU+MSXuRPs8i0/2+wScToO1h8luxPyuiOoS+ZimaaFOTno1YSg8nHGSxsttEokML3Nyo7syP
ETNOeO+J0hbIAhy8Mxn/2/BxPbPL9u+v3DcQH7QmWtTeJ8NAYjcqnVbdeNdAsZafhJ2Tw+QDPiYD
TluyghsozlHNH6gsUlTpTMd8GfLL0jqxnTOMtA1bbmxuv4Pu3xhyhbK3SfVynbtAS4TABIYdBPmS
lcB+gYKJj/bmk/o4SpR739Az3CNjgiU1iCtv98k+UtDqdw4xyiu2g2KyK9jxAMZUK0TalluzeoGW
ozCqZfGs+hl5bNTDx6bL1F6hRo0DRHJTYuO8zh7UY7BzHIsSKUEe+SU1pT2RK1eksTml8bYgsl6G
6vno1ayOf4tZjz1SyzvIMdsokbZcP98nYJufPAuTrjBtx9iaediY0muI3d4FkDKZa0jrsubCeMya
e+Uo87UvPr8k5ppdUuOE7Ix/e/KL0XCEcp+kcdymUVQht7WAxgDPXr58TthfA5doxMbliibqEQCT
T30LmtsZfZBZhtbW/zwESFY36qAEu/4AetFUyOZY7+sg3DPvy2vkv8VZ7x8SoDpyesSkWNa9qhBY
Ywy4PVYdBpdGfeT3p1gpTZD4ZgFQ78ScokxT5P5WIk5pMyjli6VVjHkSEmSTZWw8wlrL1gFj0izH
/WoKOcDz9o2enug8Ev9eS1CsI1V44bSQ4TY1QG/XZyz8eEEm7z7nQV9PbQ9IVTm2s1iVC4WNn2hN
/aRnli/Ps4//8VZniMM7f1m6j8TPLWL0pyacS/z3aXOK/3EMSUiV72XJziS10gk4idVzqJ1B1Zfd
pMYXoqcCVBVcu5v+yMKTvA+4IxB3hXIaaMkA6C200uzuQzmIIk8FhhVmdmB3/wCl7YrPb+iPl4kb
kEch6/hYTlM+MTK97Zpsv3gSo7wjq01zPR0aJPN+QldmkwVJucyopz7dTMTbZnbF16te0pJcFuLp
afy7sjaJYEZVKzgSFBDM2Nn1Wq8bUP/Bwu0Vzuzt3k851cuXkboAnfBUiRUf0b3CrUUU5c1YBqYw
GLf5hSSctCMlpweOK7CzqMkpJ9HQP3/zWBvIbPoKlStnbbcauf30M0GoYYzishz9HY7+6qwErEG7
gajeppr+mfuSih30kw2WzL2a7w0B+2+NcAx4IerzXk680PW+V1PvgSrIRI3B2TLE0qpSdCYA0sF1
U5LFaPMvi1aHtyvvku/P1GpuFVQSxukq4DcSm5nNCXKlmOjsFN0Ctol4ZXOo34szEi17Id5SFZfS
wHg68brb4x0w19itA6Fh2h8cZeYwh1f4ZJC9SO/pSkQCza1x9TdSTeP9Hs+GEX2mFJKdzRhWmG6P
CMKl4wLxIT2EpR6VGVjwT01JG8Dbkl7M2BDPR5JAh08H95VMO9L8ngEWEWw4gmwk82JJ+KmmO73p
GI7+PbTKlS9Bn41d1Yb851US88kW7IndhOSO0/GkeuVsusXmBXjCnR8Aw10LBFhZAsFRq++E4axM
uGZsrA0oYlw/bAD1D5QkaDerkuaW+DzvQ2QmzBKrjBlm7RpeOwZlv1eJVp4P9d8ANuKEdcNEm9VF
Cym9FG3oIdsrunj3OICqoWTzDEwoQd/n6SPDKMzpGyFE8JgWQp0b/Y4Rdrz7uH5U+kuJaUbLE10o
WBJOJHAiCpNteXWVG2rd2XwGICU3wpKaBoUtq7IqYpPWaa7kPGKSWvTDIVvAV9021rocZ7B6KUg3
AVNjZM+fgdvg/bZsZN4v84sMszn2E7kA1ltn7htjndiDHANM2j4yVR4e/a4U0piOryafpoQJL/a0
zZqYgaRJa0jpY5R551NOBEmmswB4HEqoi1ylYBvONyoKASxjkuL2Txj2IchGsfq0VG5qj6Vf8nXQ
zWZgdHs//MNsNGbCN4/JuBpZXhVu6kmef+qcx9nrlB02d7uSLGTx4dCtr4sbWQGJ877pIqlDA8Op
QXmE7UiYVW6mPHEKjR9r6S1VPn9Ad/ofPBcYVnDA9WsAmuK99y3Uu37fUNsQxKYzBm299PBZeF36
dZEt4pnh5Mvx+VHbCJlE6Vt64SFsIXFvSfNPhML/vkw5C85O/fJPuybO0amp5mI8RgX0VbeKCuBx
FR15oEIcece5+s2ITA854ObxWxYBVtdtCHDNlXMUGZ8nK4jq/hH/aYQlnu/xfl6Ckqxmq+CtbChr
xlWZVUlGuGO6qD/Rb9fORs9L+pFZpt6UPF0O1rD2JLrviWxmaZO6d6I3s7gohal1gEuhq3K+/aqd
h31xfWj2Hv7yx/h5SXu4hBzI8DE/Ch5AUkdyBmxLJ10Y+k6zNhOeGExpkw1N0vdTNmhI0w/Zai9a
Jo20TPzR8VDVGByAVHiZCzKDKoWPUAe8mnurwYDpFLZ2A4aXqYuIvUJb/BaI8IJXGVeIdv7kpJ72
6KORUj22EJ+SVjbvInad7p+2Bt9vmVhTw+Cwp4FnswtRvOi/X9dIBd2n2XetiLiY65EBi2/jChrn
a2E07eFqaTTOTovgImb+f74P6zkpqGeGIboiLUJWjRUXTiLW/ON6/jM+QRiwz7Nh/A01YL/JuhpB
q2GAefXRp9/seTsecRjW8BfOKkCGT85+F7lUysHEsWrDDJT6JaXbtd5+ozRxzJYhIwUo81cfZw/b
pftbQrU35HMMBJ3cJgLCNCRWuvfAeFTT0ylVVDQ05tJv/zMjP43gXKXO6toSSSWdBBP2zILaNIRH
IZeXshYvzqFOQJgn1pJU434K5/STuBrgg5ZYCrl8xrEc1z0teCRZZBb1F4NoKVhYkUIF18abhkPo
JQj0yXrPxo5oecfWfG00izVDXdOJl9cwICCD9xbLKlcI+thafj140y+oAHQPQ2XDHkw6wRooZpHl
gtH1HpTasdmOAoquZZy6kwVB1fS+FMcuL01QZu8AV56hp0sZFZqwQDdOsJWXq6yt5jpCWhvZblIA
p3Bg86L14Jc9V2VKun+K+hUVOs6kd9pYTKN9t7ZlwpJ/1Wd2wMWZ6eJfkcd+uHUOnQklkyyUgqb1
5yoTns1+JwajeFUSqDW/I8Qif05BXf0NbwVoCCwxCPc4kIWmiDtUoAgvSDGYDXc2/chtm+YmABK7
e17OxUTU59bVgMWWDaPEeK9yIQ5a9VgHPpAuovDx/f0ELkp/xIHTKltmnroBXZsqQ57XvBKBb1GP
bUZiRKHWpDgfOe1bDufkP5Sgzj7OznRqzQEwqOEXBXtfeiOYBqiifqcW4zC1Fi0tidJHLfg7dYH8
B9lbWuYwpVN42CEQ/FfUmAg0Xb/yvlbKijESAyd9lwTY/hj9ynJJ1zAXBAk1mEkiVNfr7KXUQr6K
i+wlrkMMqvjWlObrfhM6r9AhqbKfliXmH6XXI0ydB5AXU1m+3I31EmN36Xtxv7J29gLURDG0/94X
P9Vro3gOhPQ5uBenpymYbfXmjLpzBu9j0PupH6rCDFIHRaoocoHG13FwmLJU0EPlegHod1aVupft
nKR89ZA7g2t5UonAiQ76OQLzy4xNfuYac6KtzFFc1GCIiNcx+7BnPgc5NGTqdV+RKZ6eWfl9gPXY
MWn8ZfjOQUAkpOt3pvcXY2+EhfDWlTx6KxGyMqAJ9IoRU96jdoemO+3rk9Lhj7u5135pz8Kl5CnN
IdVxwUO+uNuCPp9DjKRZCG9CdjahtyrRuDH8EqloWnGXUbD04tf6K09CMP2F6KGUQUypHZvAfTvJ
umsF1dOEAaCyAqUkGkCiL4gFUgH7wUvVAKCbCSahyyLLBaCgUr/pGZJY00yN7x7Y4LMg4a8LwWGG
0FfH9u6dy0P0G5cMXpVSlp7cwX8nocSVUHlZGdNzr8/dgtF18LI2OB7nLa+Mb7N4a/Fc6dxaWv8p
u5X1JvuTbbNdL4M++POCP4F/RMcZUCiTVJYMGgg1UlEdFQ7ju6UvZYgiJv6mHu1nJAVmUoaXsh44
q4X7UTUxWSlbngYLoCvJpz/f7Nvz4GvvlZ4rQGUtxSeYxLNpSpwDyo2adGhyq71YkvV9PV8Dp9rN
m3WdPzgUwtWW1Tfq7g4gIUwMg+t6rbf5jqYRChlzIRA0Cy0XWxV5S/flKWTWF9BVzjsL5CAh98t4
tW45c2YI8u+BHlA0tnYk+RdioDZFTHxaoJIKB3Fa9PKA/J057U2Zol8bZ6EunV24C2a2gsTMFhbw
b7ya2NtPwUSsSBjuW7WOAuwlVS8jdUKMsJeDZO426rER3CCuaZHWlKBXdB2YJZiMnT9N5VI2EUwC
r7GxXsDcY9munyZd6JEt6ARP6mVsFm1f9gPnx3Ek00wiTrPndqboDQZuTR0Nu+UxxnqqMIwFjamW
Gg5ZERH/tEBZSG/XV0yhWqYsIlyhPRKOzkTOo/Jgct8+qvOwOHXH2gr9S46z63z1grD0z9DlKSH2
OK+L8UDwVCdWB2u8lGg6+JmZ8FUYOx0Ft31cZ5qRL0f2UBv6PIMHxHVbnS2Z8NSdOc0BWtU7OI0+
EOvzmOYksY3vLEnVQDxaRWAY0igXR7EiKoXATTXJlZj5U9F5bRVuzItrR0GFCs98Z2a9Uyvr2ZAq
sCBRY4PhfStdes8fJYCGI77OAF8wuALfOO1scEBIkrRn9R0HHFMsRaVBZfquUlAkWX4EwysWtMIK
opbMPM2vYlo+Y/3l0YWZvq6I6nedrr3aDS3/e63pK9l49/5luFJlYlnVk0geDY/gM0/Irrs6hPE7
nToQlsSDymVk274z0ZLhRoQgdWlsXNSfrBDHDx4mG5dl5NakaYrESmdOxe+wZND3Ps1tSvpPNaG1
UfBDFudFMwmjRDoU/R8XUAp7sFuMQhoJEQcNVYPH+78dOStQFucDg2cxH7FoFk5ioAnPI3kVvYxu
NTRbZUe3kVMAUpYbwmAWMKNnbXJ8bdR8c6uiSX71tWFnVPrLPNN0xB6atqVxuQV06LOpUVAhOt/P
mAD3E0jtyrFBE3GXjR5+DXJmjr3iJqoBX+j2OExSO0R+sD+6u8/AmKoCpKy5/Ule74/SzkIO/bli
aDVG/+DV0CcZT1rgsx0GVoeGHxYzMLuYK+VQ7wVno3VkWOEPbyPEwdu+3jZB8o+ZVFugdc8n0KdJ
Zu+43jgPSWv2qPnjDhNtvae0qPzYcRKNUsRsi6iNf1sGolOIXiG4e2BEfP8g7+avER4p+1xHRwyF
q+LrLMoEoos5iyEfBeaULT8EIcLxZPlWlhE6t+f4SKJ/LzJNPaGQO2nxSq7Bv8+wEvmnFoJEYOk6
oDWukow4EkqwXe+/F1lSdX1CaRmNBSb0/8R8j+vhT9yL5yrRsm1OjQ3tH5ZCSSRTnov8CUz1G+dp
TeEVT9tX8Hm/lJR0SqyA1lPQ91gTG+BQKfw54qsm4xtY9g99ca/gknwxGPVEHm7r5FZyVrjKJFOb
Jy8Ms730GKvgofS9lJ4/SqXvPcJbRrXkXCq9KAq6nRY5EJ+U9Es+YprkSCV6Ob1/5rRPi8IDuA7U
wof9+we+1L5uNnK9/dAcw7zGzhvv9CHkXv9+5oky5G6+0aT5N6rcgDPL2OKVDBXsWdFFBZIe9VGG
RtFS0OVcDoWGhO3fViSVuE1/3sbRngu46Z9Ix9RnRXUi+vc0ZZo28IAVzNIJr8XwbUFrJ6sGt8Tv
mm511LXjjJ7O06BUsH+w9P2K1+LHJNQxgqmYiOjDLuAmL/4zmMVfBjESFa9lBkgpKVdAykfIITkS
Ym7oXQH+VkkbPvr8O6mx0v0nWn3A8y3Eu2P4OR0ZYRRZc6ezrxWNw5YJI/MgOGVWRbI0GwS8hpQm
qjyyysWZAVOJyK81nAb/jWz4qPZG6TYfq8wJfyyRtgqPbv4IAf0xxtww+ef0QOLr1IQhaMOwEDWq
pR1LfXS6gKxhwcypR9E5UzCnA47Jhqo4dabfdDYXqsKbVkf64BRGYJuHOa1aqfYxYJ7tr9nyJ8/c
7Ah6AgwlqMkVpVfR4i/OM39GTGuLic4Xm0o+RolQu9Cl/Bcav/P1NhjYuAeMlphtQ4JbCWvYZmpU
T+IKWl/MZn1XnDHdkWXiYF8SH53cjKxeKU4vdkQ10TYQFKjf2PeaNz1Z8auu5NOhBayZ3gzUhRZJ
QkdPtCiDb//Jq5i1feGdQIu0oIbzwGbhVIr+OEqjH6LryFIoHdpUfq2UzOHG2kXgiluMduwiwt4u
Cr8V+iWougHtmLm1LXuOD7KE+1g9ww6vuGX1g5eJWNM+X2hyGT3wbAPNys94fiL31eMORbSkqXoC
8v0Gx7N8RruOwYPEtWcR/V4c+kPEUl9dtgGrw1fykgvdP6+z9TJu33Az8RyWZbfZmi01x/rHKiiG
kHXW5Rlng2XxIpZmtb8moF0a+gaXFNXAxLcAZnz6F+kVgvicrNlZEenLxVDw7rc/IwD7ysgCFUt2
S4mrtKluUzrlJB8mxxYp2EDQAMOTRC/QR+NUkrluOT0lH+yUXowhX7XQaD/BMGC3w39gNuLDKrnP
4SOSAaiEwzjtk+rsOKdMpRt7UT0Q8BJv/xWBdWDeUCURVrQGyTHyxdG8i4IcZeDhAT2RVKZMCHle
VY9rVKG+BEVJl7WrhXBrmnm8T17+SN9ui3dAQZIDhki/00JuvqxkA29PJasGze7NTpNZwukInO41
xjT4z4pu7DkgLU7vAKJOq4EnGi4xAHLYgKSJ+yFG1af2LJtwKeBkBtjYxYcnPmaENuh9qNS6t9EK
JEgkxYTkwhHMyJss0bvoSlEuoah7qNS21uGuLCjXFCeyeXJzhj+RIikbJEHJ7eDm4Ynhbt8Ha0q7
O/f6c8u4rWYsuqDGerlj8Yp0r8+UknjrkP68cYWGBLHbbQF8YA+rOobfDf15Sl/cY886tlq3dCmh
JMil3zI0afaHoy1ExFVj0jB/T9GXh5tHZISPQaKoObW5fVPAa/s9kMoIK1TkkmDMHNrIhjVtGOnx
VtdqWAm/IaUFns9mlBVH37htQ8Htl7M/bcUqEQ0n9o0/3giOu3jhpbdbucSH+9EqSixU4vMcQJFP
gmzRWBj0Btp+YndnCHH+WHvxcIQA6jzfzllYCyWnYi8U7+lQDOknsdalF7jvO+F24pvAWa9YKEWV
A4am65zdFp9DyHf+Sa0fPZ4k/P8cZHuXZrTWmv/vLdUPHxua+rcovCog50TAVr/g6DPxM3v6k1KS
FAArXCNmTuWrl9WaA8REBZMB9TBYj6e4pnbIBzfmpwNYaTGJtp0eUVDH3glwW65M0uZHoPctcGfs
n49oRF5f/CpeqT04Q++MTiemb0LysC1HoDgewSZ9xgWhepoelcoMzJAwxGMOdcpPLn8YBB/xhYwC
PHnbGcYvY6lVChveSTsGaxn+2VWUlD2RdrIZvrOCsQWBqRl/A1L0AohhtB/zr9RMbEwu1PUJQXF3
wniTcXgJIo5qyqpY4LjJJhxxIxd2xNVMbrwWQKaWzKtPuDUosW5BI7O/vmshoOgvGf7nhbvjngcc
aP4msE3EAi+WMr4qGHMk+rr6sYep0ezOU6wXAQEi69/vcsJsQbQBBUFYG1hyJMcAxGw9o024fV3H
1IupnWqJc/lQMTxl5t+vMNoTF5837shsxLaGZDSgmUV54kcgzXCwO6krLZ1CxbQMt8vLVmU7E9Ke
eul3hRyv/s96UTLUv0AKwyqlJn6R6rXvD8vzDksC6BoB/00AKpKmWEzWJ2P6cr7XKwmKiAvedxmV
vxgm6s6YQc5Zw1Ocy+u0JZRVi0FsIog3cKODFnfKN73QodA2BrFxITrOUiRfrpogd1OmEW8e2VgG
RLjEkRan6qCfL/M56k2IThu7kV8pQPcE5VY8PodfjTWoVadTTzG47BYFh1vmVtQuW/i0e2Vmjra8
+wWOH7hPGuDDUlczSQTF+e/uwrLbFZipJ2boQuvgS/gPDONnfaZACv2CCvWjvXpg80d1rTrCKFq0
szR2M/ZPvKhQ4972qok+p9n0zkCGBJ4SmfhcZpxXqpFXfmDPJN5NZsmtjOwx52O+Zw3apAypWlni
B+xDUMdLD7558Qp3H7PaAvJjWlgNWsOv7hUjIpzlYLSGFzFRsrg+D82SQ1MhSF3O+ESQo2+OSYag
NJh7PFbfrHn8FE8Z9DpZtScuRKuR/xk2KTpuSMkJH8eu1QBMeoOzpvItK12F/AqA6HwoS1PS8Tbl
Qpqo5g2pl9lzsrBVIOYmJ12R/mSeM1Z7FaSPRmaXnOOjnxuNibjLXazfXjSjh+YMaTNlN1/kgHsa
CAPdJvYZXXmduy/adVK+55aSb/V4jaHNmRrvQUc2fPssA8AhWT45n8dPDnQpCcso5dXKH7uFc/sh
/P6z6HX0nUctURvKMNOrvAVuomkVZwF5oT52aRWpG94x3gNX1Dks38vHNYxfJ5lH9oZpmpdEiJoO
zt/rUPiEyMdDNM2H47pRjwkKM89i7h5n+2qJzqRfvKE0cymWuqLOiCFiaX/90WrPqJzjEOyrSTQI
7dR7yhITUyc1VU9rDItn29vfcsoqNBIber2n5M16L7Jw/rc+cQl3yZ8W14YVeBSQZByerjusSDhA
K7QjI3r66LsJbUrf/6rfPdqgt+boR0335QnvSyPh3sDThsTKnD8vDEY7Zh4RWSPIA5T+7FRBg0IX
Ek0heXQR1twofsc7Sc6Ti6qHA/k9Np+X9BDkVKHAHmNfYAXo0lLtjLbvtm50eUbS8djq8wKgyMCK
DtFAyrlNAHl37ped5ipraAwmkzF0MIHC+6Tg+HIucXEpT4iT71lrBrO42UPbTUYdFhvRP2zP0ckg
gM6/JFa/qIx9p78WuRzGFJdO6tmT8Z2ZJKnOOxZ5XPRphpH9j3S8DM5x8YQpXCLC//zrg0U0DzYZ
RXj248WAtTAdalW3nuentl2nWh+Xl4lJUQWBXJXH9qe5G8BFgWtOHb8f5DqEcAigtNwHy5vOUvV1
BQVtAH3tLMX9Y+61TZ1kjw7U0gP7TmzTxNGbMmybyG6c4+GhKgqlVdFlV7SXdOMkEivCaZPyLXSW
M8sbYGXpoBSRq69mCJIUy/PliFi2y9KHEn9K4NTCZkq2oVKj2R8HfzvZuY6xSINUEJr1XqHTbxp/
BYN0qfwnWrt3V8xJZnnykaU/ihjyWwxGHqsfeBpbnbcXs94SRdqbqcG5RXScfHUXF+DUIM2uyUST
dJr0tqcypJavFPxUDHeiWKyT9uzy09nRg0YPmHPWZA4d4sjvc6IUmLh9aCqm24rJiI22XmLC9TST
itZ7LaBDWH1gM3yBmNlM6In4sOKphJ/UAVgIG4KEajJbJAL28J6H/BJPHUSVWtN6MruD5MLr39EF
TM0BkeZLZKBET8RNliZSFoQmbBA9N6+8DMyrnH3Y2vNcUAQ5o9n1TgPzFUeG49Mw8A4j8GRH3taI
QASjY4oKtkkYvPJcFB+sCKoPqcrAW4osi9/rL7e1IRm0cxVxxfrZvOu6XYM7x8hD28tknExdlfHH
3anZoZ1emY8xnOFic+Bi79Y7xOg6ZFNsMNMu3sOWmNfKDcjslfiSZZULShXm8GVXrbiWn3xu0+u6
MJFh+EYTEsDJM6YwwyT2xjLjeYA5WrW6BrBim4ttiuDaXtu+XhAbFCVxNkJehZ6r1UD5Q7bsruBi
8NVG3aKNjDJVzILnratul2wvHy+CMQ1hClMzTeTW0ErzcPLKUZtGK3LqsFKKMqENxj+XaCduiFD3
HQVFVVDKOaZW6092hUWqOsyevnQZu0OWq8Xhy0uj/Oohz6ilbhedAm7HwICBZbf/oPQHmmovg8Iv
fn6m2XR4/uO8swHGzihMV61WqMaFOB+07iE+QEyM1ZWcbBvlJWjNTT8iYd5sFyCUF16zRNArw2gW
WRJcc/d8Q643TaRjj1hODn+M6al8EvPDV572x5yb5aEo9gmClbpW9vqPkZlobE0oPIbRv+lrpQBr
IBOP/EcXOPl4cMvp5276jV20WuaQoHhs9V1fIxg167yBjXZ0/Q2ksJxTxLyz7QMFgIZxtpj2ImTr
wwxXCEcAq+4CwfMEhOsgM7C6g5mHcjUeZNFiChO9WlZkrudOGKcYz0Yao1FtRqKohf69RC4kMEDX
Hwlq7U4F6gJh5bWtl9UpL16iCBzwywrgXSecy8J5M18GL3tAMLg9DvG3LRgjZ3m159ClJ5XHomEy
Hs1t5NRr+3etEu9tV91zlkkcyCtnYreGGTePDGBvclHQgo+F2TWKN3S4ueKlXatgqazCfO0wN71f
9H7BtrEDz87yXRITc4GnQW6XjMOIN7Md6dj3njaB1ywZSbNK5X5p6lOWhxSZxDlV9qY8BtbX83jQ
MSPpCvq2UrjoKbnCCm5ZgaRPBfHvx270PBfkN3Q3psb6j+Mn+ICXPjiJI5w4QecGYh65/WutjskI
+76nJdnmDl+Je9GNghWq4SglQInsRgLegPuSlVJUpVRb0J/4bgGlyah4ZbILMpFGKy19XLUHB01X
vgO7Imo0NNQIw6l5FBUpOa/AG7Z4N9O1BoTZJZgqvvskl59wcMUsFpmGI4RkiJe50GNrLH4dv9Eo
QaFxnL3iY7xJpOQMANzKPGSLbC1GrUhIxWfEG8IaYJ18K4VXtdQmREgVk2sP47s7vm8OYt3RiC5F
tE4cJQQgNHspwvLR96hLCILIjh65IsBZV4x64dJfJ39N59EetPWNtF3XDo6TCd2UN/Dp9zXvR7oj
XHq7kWdigSsrWSg4r8hRAcGS8sO0ckZZYNTsbB1R6+ENe2Y0fwWuLORe6ZE3EQxhSXmd5KkbXV7F
Dseteeu56Zwsz+rxybvPFIGsk+P5BrOTRYdIRtkiWvzSrPrGWF2lPs4GniPN5jyUyJkk/XM3tzH0
/X8fUNqdpN9V4yR20UzZAQdyFKo6bJJOIsTe1hkgA9q6fv8NumKvsDThxyuPncwOECF2HZYacfry
xu0b6pllnKo+7PW4p9Kkks4jhHPzx4UWp9yJqIHU3dqbEkg0iWmNAgCYp95kQXczJawcw+6C6Ebe
PKz7GrupKul2uWdXEBKT5QT8olXqKHq1AqYQhpM6G8dY1eCqnZqaf+Cawav1csOI9zAHAdjwOYBR
U02EL6YkPJ01M4VlTvPE0rfOZ+EIZtYk1iQrASo4hElInZeeJ6O+r6hTeiP9OKvSgJR36xgsShM8
c0EiNT+EO1M/p3psQTtAemecfOUuoR4VAOGImLafIdaqZEdKtpY4Qmk6sUJO1uAvKQUyOyD/RKfH
BtoEOByuDZMtcAa4SctHEe5VAb8kNfBBvvUrKd1nQmETRE9Zogi2N64xUM+yZ2fDdIWfge+kI1mv
e8VrX69uwxNGJzdBXPkgiG6l50MWYRVNw+kirkPl6UujExqh/YBlJ4XEpcvEKvegGo25z2GmQjUC
IBg6BfC+kgMc1ygval6nizfpgI41Jr0shObzC+jyxw7qStIzeVjlczvuMQ3rxCsmrAPOfRu5I1Yh
wlJhp7vK4E9jtEL3R40+7gGHpRdJZFbQcwjwHSEu9sJztw2rMe/eoNQzsBO7jf7I4ksjjOPsixRy
30O7ChctMNSfgWEMbIZoDwyZVnyrCvXQ9LC+fjIUcrs11KEH0mQ5wg5ldZ9ADUw+cwdp97OMskhJ
mA+/R542BZ6+Ap9zFjS9N1p+XCM/CZQcufjf/2i7p0MaRZo5pWFYjhQ6YKMAKgVexeXUmVYcp0rV
eHuZHgedgrX+9r6PMlk/GLvKBUeGV3vzUP9MYm25gUIhkJar8nj7UOaq7PuwtplbvFOOVeEaz3YE
lwaa74muONWkqf3ajj8LFTJCWg6mh68X3Xt3UvLCYPEvkP3Qq+CvIqT/uaOk1zoYUN7xBw+zrc1M
o2gXsnAguUyrDpQhLrfF22eWO1D6nBv+w37scs3Sef7tJSVYM3BKJM+mTvl6KX6OXc3BnvEMSSXq
iIfCQHs/A7uX3Ke5sEEjjbocN11h1WSN8/5bpCy8nruBif5kVevOY+lC7+6saJeCUIjeKp8Abe3V
F+JyDrLIZsZqEw8KL+DQN4824opKWwQpFWzioIyfHOL+sRhszKly7OAT7ndFv1Eg/bjt4vUuTOBZ
z+PxvJn77OeFAxjKf7ZshtsDSkjW6AWobQalFhmGIQBaxqiOBMy+RkVsY8gekn8NRnykg1cbq/UR
0Vuh1vPBpKvqyOiKhHsyEYLY2Or+KF8LZvNZsvGLa+afSRUxn+S3+N8sdpoWujpWIxdvAOyhhu+2
u3B81xXKEMq8fU5ZUeEl7idGj5ttgyNSgPpVr5V0Wl/SijYQdoa4tZFDi4FKyDymZUQZ9C9UQHaH
L9dO0sf16sjS7ehuX7/c8Ob52uqcPPHrArEZtZNQjuNnCiIKtdDM8rPDdotd1S3myk2SsmuDyNDa
UetMvz7kFQ/4KtSb57DRllNVzhVKYWTzjVohNEPJb9pikvpVY7hWjTSG4v1W4OtMfd9b7FnradNk
qAXJ3jldNxiUBqC3BBjjfqwsLv4FRRzx+YwoX23xzfqp/CT+6q25FK2HGeW6YJ8Xoqn+RZcvz+7+
aPUhfsdFt1CDeFWeuUM2097wHrK5zrqMb9TNs27wVbxwugKb9+2WcOPdHQNyE6JA0XRRTKKUfzbL
08ucbiRUt6E7yQhX6mhIyA4CH40P7D1VSxJar1y2AzgU8WXG/AWVVAqWgtjiYLguZ+3L6nwXSssS
Wzo0J6jQYzotq7c2v+f3shdgjHFlKdqtIwj6mQrqmV2vs3UO3/zNaJXgX79TvCjw0dCnxOfvQa4t
n/LayW3rVo8tIBwkRPEXemq1HzpSRXA1gIFrljGYhkRZIxBf7ezfDJ2z9zoDVaAI4RSdkBLK5m1p
0lNqq/jpQIyZMtPOMestvf6PU8XpPB7Ei21k3EbbVY8t8/q0bqODDDgrj9Uc7AQPECTfB2pUuRN/
mV1jJ/yXiwdqJ54t/0XVzVCh7TD+TSUaKlAxqibKuY8GwZ4+YoemCjzoiuDRI9aqDcnfgENIWYW/
00O7v1mojpKv39RAhkjxMQ8IGupatKurppwMRFklcbX6BZYIQMi8ON4HsOpGPGyCzVCnpeq9sgaF
OoAiJ27FqvExnCVfEM4On2H042V1ocZZ8dG6/Q0kcIiFYGWFdeWFY5JYOcKZ+XO4zKAPcgpAKKzi
anQAvuEH9gQO4qumYxM9ixA0E/KlUsrteK9X+fVotBFoctfCbNFV8C/vB/Ibfen/ZbWuAoNfQ9Ym
CDfsyenFOQYth0Oe5skSL5bTNOL1sdMn07JKaMjFsKUBJw635W3KMpFk9TW9vq4EeEzy9+1lrZJC
DF5IpcjnSvki0ki8YTWFL1f/3PTkTFGxexCgijXgpzznmwX6B5kk3zzEe8nwHRvgL7vk2vnFVmsl
1EbqM8UjjP3ZE5c61pD126f+o7E2L3jUH3Uu0AlHyEoSS0d1h8Yi9mJ1nxc8PxCuktI5uhT8o9xv
zPBu3CHwWQpGm/kvpfZecSYjYgPAD16xIcYzU2qAZmLAVDyPFRVr7BhvrolkbWWg6iXNn8xu38Kj
QOPA9zIss0lcUHpNZQMcs0J4QbhVOuEvn5eNKZJKWlSi4Is43j5U2CZh1X6oUzvHcCbfWBVbXt+N
f/6jk9yHQk4RHJI9wjstc2oV++PMm6Un8c1tHgLH+DEKBtTy4DgDmYFYYQVmVlFOP8s2IlvHZqmy
wSG8SDuIY51Cm+qr9oAcin+2QAj+6wlzCt8/8/jiXzRCY8Vhoqon4Z3ICWSagjGXIiuPRivfrtj6
hEnf/p9SFnASfbYg0w0Ph5Im4qrzn+WIumRe8ccuqh8v8K3ZrR2ePLcp/iI91Dr5Up4F6qVJYMLo
bENU9qe5h1h9rVhG9QFiVNYnQfroCB0P9EH8xGEmvmV5fbtt/Wb8OGJbO2YmZ14e1l/0t/5DXKJd
QTc74TSdsP2uF4B3I6Pk1ILcGoo0zY+iHuAQSqdZmSIN8dW9NqlqyPRcJ7mjym0CwpncVDCCa8dE
f0wbzI2hAvHY6dfNo4Qmw2d1oDPTmIaohroWfKyZAky14VrXreSJvLEyX8hpTD6R1JW3UUsCcsEK
HXE/wtTBwJEoFlxSDfPx8ApT/GaKQAZDnJtxUk6RSjekwpCK65njLa4BQFclpc9Ktehlx089trRt
2yt51xeL3Rd4NkLa3rWultP8W7J2VfzuKaRFUEn3yGE0CyvwZ5rhhW2p2nSbwgFKZxv80CYEsHFF
cgyCk323PEl8rjSwtDrixVKY5KkYocbecQS7MkCiYQjvIWQMeyKH++sAa4JjpZIBljZj4r1NuW9Y
Kr5kVojskn86XZmxW3vO+X7+X/RCHZ2j3Nulsz6Qaaxw+JqeGxT1qe0vie3toT81a8d4yGHO1IS2
USBWHnj3hZigJGNUuhRjQHsS9xyMTrOHgZ0qtu+0GuylHN1Cx1B7fC+lFHInqnUmkodR8uYLAYbd
OV8tsauyGIS96GXVthozX1psGIWMx5HhDNPRpUQW/9goccSe5PPjnKb45KIORlnVB5UakfQAvXSo
Vjw7Dji+iZp2DeUZeJbtCplB+OwlCSWeIUz3LiLM7h7AOLC+/4FwlMLkMbYzgwfhTnbxHi0+DrB2
AlhF6jB8pTKELcNtwm8XgqcA3QUgDnAPbqgmLmrtOKCTE2sPURja2ZpdHH9ZWPR5jWTbMcAlCXqf
0S1DWp/9GmZt2tU5zVaPOT09npJkmj2ZZwTYfC5brATnartjpCLUSdaU9dh046IzmuSS1hUNGgQl
4RHB9AviA+wcePAOducLNHZYjC0il3Cpllk4mmIYUkbK7qWR1tjZswwmYMrrK4BAHzOZiL2JM7d/
Pc27cmLoQtPgXq9V/8qB4XwAHx4p+R1aFnsgSKbtNjLwky3zNOZBJ5KvaFLx98m0D9Jqp9L4rWTv
+sL2e+JLXdS954Z+XWueHcjkc8GCU2MKcQNGZDza2nGJ+e7GX3L61wZ8wN8IpurLITviwEbTYANq
W6B9u9v+YaixhK+lxtJTpVr2XbS+W3/TPQRrju03F1KO3pK44v5VV/cZHMlSb/kLMljHsbE16N/k
3xoHP1bEJGYxf1q+H9FTZQuOp8cDkvmj962NkLdSzlOAb/00LC+gG5lA9jsvC6DjLBXgk8lnMotQ
1zuW7kt/OoEHEckXaFvIHeMnLDkzdBQKzNBlhqVFbQdRVouafoz+3Dtn3mh8fq5l43zX4SAfmrFZ
bKvr/T1mFlFccz0XbrgqHNW2pxcYAqg3ku7VBwWYyEjKdF5wMGA1oOrzYxABZmarJ1VFSimdFjQy
H4CsbmejuZyN3Vl2M0j7tECZ4pUXMneAs5OLzeOvpz2qDEbpxAue14akVolmNEUNOeZ173EF8UlD
FiKdE3dZo1ZFYl8eqgtZSOE9dFGAiKY+SfmUAlBIaYYYJrHqrR9+6ZNCbt0z7vZuAOwPM+K1UMth
4Pldh7nfHSnUJtVFe3Ifl9GVDwtv2WdVkYq4ET4zpabSJg2DudjSNivwjXWl4Va7y93ge+Am+4ZZ
6o649Ml0OJyADH4yEb0DPM4smNpNUb0MOMHD3MgwRaFZM/N+mi5fQzj04h0Nbxra4QFrsoju/80G
oYYXFGTJv5bKbWxYnLhM2sGRzm/xynGwYFJKXUNhj7BSa1sQOCr+11jvokJivvn7NhM+lgtn5TLj
gWZZVWbXrNX3fTDGfkzRnNXe01O/XCNJXb8QEhp00Y90gg0FcUJnjLlLYkybKcJDMhv1/jkYkjKY
uYbSSt3gsUGSYE68cWWyJjS1Ut7OlCYWoZJu1nrMOUVNX7ik9/wSU+hHCvn6xy/T4bAK0CtOQCWq
+UnClwmKk/cBj6A+2+Jm35E7FEdQ1jIsIEq91SkdfI3m/MPr/cgJKv13KKl2grzrQy8l709SOUB5
TYnGwIcMXOBktOL3KigeFFefIthkbbWlhY4G0H5kxOV0zJxEzOgQlgO/yRsKI9BXkGZwV8SauS0+
xByNQoV8hYG0c5I0M9+C+jrvmrO1ZTPBKSMI712EBXwmBcDjBGe8/1CD2z0ixbncZemSO7FH/6Oc
fhlpDy34oHdHJb//B4jxCX9KLIme7HdmputqJ6Sw6BWPSgmVFoMCouFwsr9sdlATpynt/iWJnFc7
ttjWX14SYIumHTCBq2aOCpEXjetebzUeyQ+W2XvMUf4qUToBIbkbDQA7POobXy8DDTC5rbmqXVW4
hnfKrorymYJcplJh9ZyECU8uwVDpscWPkJsIc+cnQ44cnxxn6GWpSUba1N3a0FoUQ+VkThYCEIso
qIYif1W4yuHQIzRGe3nWipHG/N+m4zchZO/kU/nQPxCLFW98KYj+f+CzG5daGVMxZ3nsywC/dDqa
+KTojLJOV7e9Jaxj0sXQiTn1qVSwuSnbYuDUmpwvl8FnlTLOWP/appcp4Tcjb7PXZWvWduwIxfVA
kOlIiQEzkoKpQK+Y/qjjbMsteJ/TOqyE2OoAbhsIUpfioRhFjIRGPWqSoxuq0clF1jNt0J8mZYqt
mgKihbsTMPWbt+F/pBhccVCDlp+MCrM4n07mBBOd7b+2WTp1jiSTmmzKYK98J+QYAFm+CPwusxEv
CqM1jV8JueuDLXE8/B2tD6qOXIHqFsCpOV1SW6AFMXcIR3BzUVuJN28QlUJnOHcGMLHViBn3M0/S
3BtkvtoJI7GQbBvbaxHaU/PD30RpgVtUUrIQJr7oVDMpq9pZZa4yCi7qDLuuhcjpODE3tZDsUuc6
f9LD2ypVPRyVXoVlLN15dPb5+XHdmeLfSup2YAI1w7W3LvQR632k8fHppYoOSnhv/CjBGdSSWeIy
7N48zRXQv/qaB77nL9L2e7oKL8OTxVHeLpcl4rcwE6LcBFwXYgrI+n//bE3XE0iXjMjf8Qx0os+g
rM5qryq5R65A4HhhigloBBZ6ERr1CbogsY3k6MmIAf6ptPs3sgUOPTHlYjqlr/0er/6m8B1ba2t/
3s2J1l3U/XsURAkpmxMsyTiqil6Zqa1ebXkXPwRUZC64jlOwYEFcTlsgErw/XWJQjoFEaxkMPEj1
NXFUe7vGf34k4gcTsdtSeXCYDdtWj04P+/f/nxOzErt0N2bkfUmcva6VJMR3U+d53sYE0MPSAjzR
ZPsJ4akuphjA3DhNgJ3whtWe0AlZolu+6AYQkuv13Fhej9EGnrUPhJFXWrhwCG5ea9mf0xZeyzYI
TFfWDgZ0SlJ/3ZHTa8qUeofxAQXE4w+tY39kbT//6cbywRsUOrv1nuCyWgTJ+tyF+R4IaMVPwtK7
qStuEemZx1NwuoDKUM1vv+rkOJIwqP+nqnuy5aft+3o1nFe7XG8903YjPSsCQD7uZKfCckycwQ37
XXT7bwjfT2APWJwQzPqVtiHSSqZLMmrzzkGLbZce/35hmJUA8HhNBH6fZdKMgX51bkOx2+uDmsQz
6WOHjm1nKYI4+ttYYoSNBIvgawiyMtz0WfBTNeWCwW3tiLjq9Vp1NioVoBcVzVcrl/SIOEQGQvhJ
uPqaBguy+fkWowvIB89Ay/8IJ9AseSWehlzsyNpvyBTBE62QuMoSql+SsXpmafb1p7HJw7TUFWRQ
EO/uHpNI7xlOHyDn/gUhUs5+1XBUnk34AejxjJq4b9sc+exqKiCl0h7YdG9KgDD/Mas8JwHBbLSv
7kXqE0o7id4GfCI6Xm7CNLYTivjIWYpEWuo5cumzHt+zYAp5romnZjyDDUC3JEX+mrd738y7D4xF
VkDDa9ZubelTSa5MB8QEfJ/ANdvZ1OOZ6NYTFHuhoWx7xqkdClISIYQpaIZItpbyFDHNuYeZtvSM
a9wrTBaXjLcSTxj2oVgnWQbHgdwHTgOFl+J4pZqKcECz/MKg7OkpvTDqCBkWbnrCBDPy9Pczm0uB
675VCxZb1MKngRmJqoLkOWhPL5YkGPUGY6yqGeelB7AqRT69PXWlzFKtSCytYJcdimws0U1Wtso2
fm/gUl8QD9uOfCgHhI442nta14/28kJp1D0FLQQ09xx65Y6Jxv+Lh3JC0+j88mcpg2eZD7YhPrCJ
03QS1qXjYOiTQrB99b1t2gDBiV4JPfguQOLW62Zxu07nlneeNDX4AHf6CmFoNhzebKY0UTIpSpO4
xKsvOs+lPgdskZmbUtNSw25F00eblzRo6pp4+/pJ404h9ypntIG6iu0ZeODbLHgMHvMxI7N0eSJU
hGAy6QxPFJctugg7z1NxKw+aAAuyXn/8/biHCJNLUS4QWdXC5trRzdE0hGax2HXDh2j+vGvQkZST
SkHQx0FXUAajY3GEBN+X3sWFqv//FdWf4XzQv7DIGzj2a6YJQ5gStcOGIZmiEReB3fPcfC7B4/f3
OxhKCoIM4Et9guKQeZs0SlMQH6ehkYsCxYnhh2YTsSt22A0rPvUGjPWoiggfYvY1e84eHy1JE9EL
hKFKxLli3Cnj9/J8OAY8Tbit0jwc1sksJP7np3/B4CgmbZ/xhztoghlqkkrPBF3LNZeOsCJNsuPI
UTg019oI2Hsm/7tj58FowqyuPmCgyZN6zg+P779yiz0QSdWxKY8UvQlE3QZCYzvsdqYf23IWhqY6
Qp5u1nemRAhwhH/zY+EV4IGgpm8sHuoZNXHW9ia2F1ULWXlW4TejAlyRTwgssCaynhtyci00at3h
f2rcnuEHmiCzHcxQkC47e2/vCImlPdyqWKtWvyYSqaVFxgAPVa+7feRJPSBkI2g71PIQVS6BD2YV
Q/uqz0WyRk4qMFWK2d8dbE5+MVs901jLZzFCOpq8bUfUt8fi2UDR2dnqFcibYSZyoKOhV9ZMcIeJ
76h9+2iOLsJ9/C4oRAckjcBU+RVOCjPZdeEl+iqjnbf79b5Qe42WZqYMhzxBjnPg4v8T6+t8AALm
8cPm7yHtb5zHZxFhenet8flXRo0BQ7raFvuLdFsknIPEY2Y3BrlseCp2gPk3ndGvz4N54niiQ4xI
FYJfdI5xxyTg3glPgLuHhAfda0upIrOdi5l1LSBM2QgCE6txl/OVcqC4o2J7o1KxoNODfJCDhOBO
BumMwSS4LVZswW0dPDVrbZLYHeQir9QZE/zbJvfSbdfQSG+7zJys79tMeYgM33Q8W7Iel/jwrFi8
GROoEkE/ABC+T0h033pkpHRpJaxkeYvtxj3m3BqLhrqaEnESsjoGwz9AbnYtxjFKtnkOAMwSaO74
+drPvR4w2ZfQy2jriQi3DhvJ7mrzThxc8kqsdF5td3uGESJeE1JdWw3UidP9Yj/coCdkHFb250ii
Km4E1F6IFI/VCraxD4tQhYNcjZIzyq/TLdTf3Thq/lL2/wttJ7qy+ddFNPZKXsjjTZWxx7IKe0oa
8n4qj7/XePruC0nolaxGBqvjE7AUinUGRXEQw01vf/jUkFlR5+oE/trkcW3vmWQkR5oLnywyoCcu
fNcJENKK3XMrXzEIb2kKVnVhgce1k8lVsdlBNUvO7Lc+4KLMpPZMPfimasvaVRx5atPHqUrqRmu7
lvjYPZGnMk0QHLH76zi1xtXxOB4OpsT1BSeIiYjhM/FdcbJvmYZT2E3JSjMXR7123zoW9BlXD15u
1g0YK5fX2toq3O0fs9fLcOgicz73Ra3HzTEO7cU5OLpS9MC8/biXfizSHMUtBzbvVmA6As4OTNDK
7G9G9XnD/q6Vbvfc1F+yDjtRX2igCV33fTaMZkmpl2v+LI0hQVDVXYOEgv12LHMH4J5KcQsydeS/
vXE0PFNB2Az12dtVlwwWoU/r8AnEvmh4mqQYyLaKRWklDqqtdP/3iXVyharR6JZbV11Pr3SJr6Q7
OEdd4nkY/uzhxCGBar+RyCwHuDN6cc6roB9s3ktKzihkbJjaSBfHnTuZps+jME2N2DyzhZk5AJNF
u4QOOP7viKGpuHyndRcZMCgvL7DRPMQdiSyhSCUaFVC1n6AyoDHNQkChGhfLsMXfKr2ywgd7Qjfw
GwmUENvhNv5awv5ALaBH9CDllkt5uIwzfXR0VtyptEGmpDQkZEmnfE8Pi1aq4w2itY+o7BEqjANO
QXAKp3M6s3wjhDeXoHYNElihGcQh9MPydPvcQ28CxgPz6RcXxkB5HZW13vywu1fTWwwBdF6yBHfF
JxAXijDbKXTqDZdZsEANctObGYoThTY5XbjWfODlMu5XyzZs8a4jbi4O5/p/nBM6Mcr2vG7pQO95
2M7qhBJeQXwW8QDAz8gVBnZerHp5MLHzdMoov4CfECBpY6x5OGmrqcCD+GJyoD/SwK1JpHcBUDcs
y94e/ptwuVpk/Weu+tj5AgHShQwoTit+M9zBWu8x69amveDVcDV7IMe9akxyBxjmedoRTbk1VGBt
IxY6lEG3/8muvhBZJF2jF6OF4MF6uqy4aRn/fX9kLmtCQENbmCcJjy9bllHMda2Hb4H/8uLnf2Ok
C6ha+GL4xEi4xF3x5Hbyzo/V9ZgKB3G+15douF1iMlusWzKiGDqkvXl4JJfBamx4KUxytA4W90IN
IMuwj+OS1cHn7NwBiy7StVaW1jLNfghCWcmxiGW30iNuvFmuhU8TXNI+ICW/Aar9hNJnR92Dg+O3
ZkiG+h+0ttSoQ/yAf8Npzk6aHG3jW4aS/GBpaRwqgKe0RKrweB4LsUNJ1274k0NjYRN/xJNuAK73
O5BQNN7gmeAwS0JGJc8AZGPTiUPXRp6Iq3l6ad7obOcrWpJm0/80N41sq/Q4Jo5IjOoOq1+3vylB
w3E0ouvoXM/rmAHrMGuTZ8yO/J+aOhIvG+t05DYFCr3r0KiBJ7gwP6KRQPmlJl3/8LGrl3E8M/Mz
IUWA5z8GGXV8mx908rcBdSvpOUPubnrltLUeoQw4LF83CXsFj+PXDH+ahA9RsKcdkfH4Fl8vaDbX
DKq9n7n+m60a1nYS5KaIXqhTSAMZy/+MQ+ZrIqQ/T96QZGAjPrGSRBpEVDTdYWCkKrtdM+CRx1jo
bPSbeboIItXBrsNFFAFjBsYJm0dJO8DY0932N5XwyDcpubd6warslxRiwg1l+dCDySaKpWH14pza
n56CmRqroKqrCqMOcPhcwFi7jCOsx5Cr3tGr13WNe9P6uuhp2ib+vFjiZ/Y8mnUSQotNF6BjZ89W
uP1M0Db//j7soID9cd2LT74rrwstktsLF3+7rrwVABgTpx+ewa4/2J5W2pA0tzBZemaLUbPDBG1m
mkFVynivfX5L8FGPJ4l5knLnwTafxrxL9tgx1DsXOnk6MeJER73hXwPuSON5PNzTnDj/HrkQybV6
CJo1p/ClMvpQIwIeJwZqynaLo08sUeIJmRX/5EDSbk9NIQzU1jE95a1F6uWKl6b7jPlaBp9f5Cnf
XVwp2g718QNpkbSOpLH62xHQ6wI6sciAM/j9tAf4jh5Rs53LpN4+KK+Qw9xTs1rAkl7IQH6mKMuh
RtK0xWdxCzKDGMhVSmZnAQgAeVmqGNUo1FGH5xKOEkcqUCaIDh6uSnjdxTSQG+fX/cUh8hUL9osn
SCbdpJ53qP8rO9IPWMzSprXUckqkWWOsJLIg0TtUFDZTm6iCnSG8bx/RXDw9ToaCQqOIU6JXhbrD
O0l69WvxQ8/gDNzbp/kRjQLrhgij/WIfE+SpwvUT0ZWky6cDtG6zMy3tGZSGNlO+/m8LkpJ1XBVV
n2N4YdR+bJ3utTNK+yvIbg2moUSK8EuuX7n5ODJeYa4ZYM5HqqtB9oBLN7EEzTbZIkg0A3ABfip1
tzI/jcAv7ZygJi3SCpDTsxw4HL5dZIin2vhHsf4VquhFTEWS1lvQd0TwkTkxmcWX2rkOar5jZsNH
LXvGVCig/IwJn7+d32UYBBYs173o4prvg80z+lNLM6X1BxjgaiO4KDEYt1bK2vo0etEfaLv5xCmY
p2cWNssZGGisK8DShiWwQmpICroczZsoxxt2zz0d0DNSgS/6gtLyPyjVYWJrk+r+tZDkQ0q0Abud
OywMLMre/VXloo+BLLq4uUojOAc/aw6Zcr3liTul0dfUpDzDnKcfn2fojpH2R4w4RUadcuUI94Uu
kFAFL/C29D3vuZzS4H3HKheOWno+cqVCA1DsRMK8ljU91sRrCp1P/2ADhVYiqAmJVkswb9LmFQf7
ZWrcyCbPVvY9H0tyBoKHEesHeUEys7zFt+Ymu3lObQM6KWHlLcDozayQEJnddpeXQ+/xtJHRsnpW
45eSSqx/awBTk5gaGzZvclJ8yMHD2Uhh1GuEiJvlVQfItK+zZMQROVvDCf0noNTfL4O2vEkv0Ihl
zffROBHAcRQoE4Mcn6mEVBeKRy4MCAG+34QukMWxaBAm+npWk57H8Lcc33WSRwIyvAgAg+w7eqfK
NaIVEmTOFwZdCGy5TA38I3WZgY65Zz6PwF1ilDELEFSbMe1ttyrSXEeFPgcmX1lzEt7TQSvBMNi4
IPngehMG1+s0WTrnYA7sBxYtkKqp/jU4Dcw73QLx7wyRc7+myB7iJy/0Zparrc9W1zCV70+/VMDp
Va3IGGGjrMfCnXvosIqv52eyueNRC/3HrUrfuiGBlG+RcYXM45SSQYO71UBGEl2folopTx3bmcw+
6C3yS0YVUcxtfJGd3LTmerIAqqiJGSvIogkDviExaKfqVZjwIvrav5p8u6kTcQ3gfEBf4R+BA+uZ
lf6WMH7maEXq9Xx3SlsIOnuT44VfgrHMRraJ5kV326HPjxeKKtAbneWSvWv8091OSASaA4ifjGFJ
0D3DMAmuoUxDE4nBL+X/5d8mL57P6nME0B/lirIus2CpPBEGx77jY7s0qrFzSd1D50N64dvcqRhS
2NKuSGBdlrqozyxR5ldz++eNG9xnqx3XMpi7e6GAgFIfSQVm3YURfwTe6u7pPHp4LOZZhfpHkAPB
/hmVh7mWXGWE28bRwi2IaGpll4oxpICDQW6OblcxxsNaZ5cG3BA8w+qwkkhB63K3BMpTySN0RPLP
THen8Dg5cp5seXoOLZ1YmDEMx+hrpGwhAWM4DZUqf5YncyXdtfjwp2mMVyyc0CsBDa7dfiiz52En
xGVdUK+GhO13tupEMAFC3E66av92N7VxPG5EfGceMiOTgOLRFtq/wd6fSqdUvtxvc4nbC9JpPD1f
NjGgGr3SE9YhyGWPKsdBJT8wyVimfxS3/hCmgTSctAI5cR2ztEndMNzfFO6UGU97/FCD4SDHp+a/
jX8ajcXvtJK4023FjyW/OiAcKR1zM1jThOHEkD6lciL+7EUP4obkm9dedExDTtrjI42iIPBoDddU
72em0RTQiVyQ3dljxyelvg4tkG5qpuyjGcbXuoHpTjHko7fYNdL6aELRe9ZQG4k4PYTw7EzyPLg6
Q312UKOG7ud+sfPgXf/5PfmurptpL156VRSKk0+zZPwzDClCU0vEgD53PgO8snmct3jKx7CXNDws
g2VrceEjsQyoG0hyX0B+75CVyGIP2SKxf36lJ4e1reMbhc7nw3PTNY/cZ+j1kIFF/9solLp35Uvx
EwAFiwRjhiUya+Pkz7InHWC9mO9bEchENVSxg9vYw8QgoizpurOq8EhF7XD8q8f+khrc8HB5IRcZ
THzvAAGkMTb6nJkVVLREXjrJ5cXOWJimRVAdAXWDVIZNMxVroGtNssupkDG/vVB5JOfDcEuLCNr7
QAj4XTZj+vriw2cKZFIUhSdGyTSn64iOFoesN3yrzI4/21xTzi9Cu9u0ij/y5bsVNlFNsKoEboZl
Tcx/wUigMr2C2DU1z0g6oW7RAQ8R3bJH/Vf9noKQWg6HRMoeIBRSjrWmaAoNmZJSuwhTdy9KF5+b
2+D8iD3im6g8hgBf/6Y2RDNmyUNkuO59eZo/d/fK/Pwm33sIQ3TdgvXH+IXgUKDeH3EURC4ldWy4
1PmZtxTzLT+9jRMHO2obS2F7/w/NSEBLBeVGqrRGxKD2uYSIGpe9MDiDL/PUUdKivXoQ+9WjPWRF
0mXqnzoXFOPxPxysez5z6S6iFiSvO5udwDnqIAlEeVp1m68GWrOegw5rl0j+WZeHXjOlDE2vi+si
dg+JnUin+OEILRy2Ts0F5MWNNcE11ThoFHxIXjks7uFG3ACIhi89ki388YeS6kjGY5tmFFuGncOo
JLgynxa6MEcoyYyJGB/Kw6ZbW7A8/RO4D7WDEo6hYcuNPtxbCq1DAl4Kgle8I7d53RvUGDh+BLJ/
rXbUqFdA6FjqkrGdCMqh5IiGC/64WIxj51WYppg+1c0qlegEMFV87meROPF+Cxvphy73CLCI/OX7
etz5GYmFCXlF/GAE+HJhrQD6Txtd8xxJcfIsngnA/o2Vjwn7E4x4Yex3xsN+36OgudpF9fupExOG
zjzxGLmb0hFTPJ/WTZ5+aOkPUZgLMql+VXtGNI4YJxjTa0gDXuWfbz2mw317Jri0k1cL7UcLHdT0
+kg+szwzQf16G9l38jdncOFEgcy341kGVasS5wjpKqyfa8pwLixYqSkBMFkLVgVY0uX8y+S9fKay
d+OThQnL7KkR6UlgNWanrvNOmVSs2Y4Q/6zlMD97jpxRbcmpjqGt5tP5Q2+oIv36IclYfjYNqP1p
IjerZDiGvlh2BLQSU+sNTyGHjuuAowNyuNNbUB6OIHbdH9723/1m3rUGchXMllGzAoge8oxF21d4
hCWvWViclrgxdg+puikKu79DmPKJbQ85WMAopRxiHNeyi/vqzf9n9Ddf/LJa8FngxEHVJdZnlTUl
D6NtbpX6kxY2xeP64ViSt4gNoAY+ApTVWCJCMrMHrF19WV2abuPNcEX8/MCuNjqyTIBkjHlN+vSj
qmOjAVtekCAzmt98/cZhgQI2/AnbbvKH/6abv/GZ0uV5TadCiwszgljyA33nAvhPqgVEepBp+WYi
k6q/+dNAJA95d2oWGF6OM8TENxOK9oi9WhN/YU2T92ZDl5tmbT/n3DyNdgWGeIyXbFEidGjs0Q0m
MKoWJRDl835s50PmlZyhcYFNeUIzj0CdCflv9k0pshXJPyeEWyYdIxtyFQyKXqWtaNFjjnqni6xY
85o1NJUpYGnvJpm/ohYkhTCrWH+hgL8Mi/MA9YX3MVuxOTHHsilCb8LRJhW5fe9JVmRRt/l3iZO+
yJfRxkrkPqeOmOaRuHrf4iQTk7tLelLXIU/7sdg4hO52882bDxIxqrI18vPb2g16hVtFMuPsZ6uM
DFweWpQT+v8OhArlCMdtBX4teaSum91mSlHTmYXCcUr9r8cUb9veu0T62LZ0ooKTXV9SgNlHhkdw
CbmDoJHLt79Dqo9RspJU51TtQ0OTe/uR/lbetwxYhIcobYNiQQrcwzJSmj+757eY8j3sVJA62Dfl
Yt4IcHOHBoF5c2WWg4uh9PIAHewWrQS2+5DolusOIQwS3/IDzoDqHd6DWs6uMgA6IevqSxATa5Or
6uCcVayeoqCPIRCS8TciCOaWshhu/f7PhRWJkDebBBzLWK8p8xiiOX1dphhXM/i5qOikUzW5HEaQ
NbbmeCvpUBPK4ELL11onrl+tVVT/3ffvSYvl5YDN5fkQ3bruglpUWuBn1Rzu+13xjL3a7RySEc+V
SXEaCsa9N0e8O8seZ3YjT0OJGU/MfvmIMtIOaG1StcLYOtPz5Q43yVHGcKaMvzq7MTTYTq4YnPrG
J9C4e+yOKFAWZUSpnHn2Mox3Vadc6dV56ZXhKEmxvB8vLNZmycjdjmaaLbyWjfHmgHpJ01HIbF7M
CSniESy4u2QP5Qa1MNacGAmsZQ8uWkkr71YEZTJ18PLahEOC0QsuvDp1ibBmfnD8A+udVPNmLc/U
j8PKBk4lWMBLF7TpWEvu4iiiuYa7aOtroZODhEfaEV6oOOK5DigYTUQhQ96CK0GM3HU5kdPXD7Vs
e2Px/+G31Kyj/0p/uazFI8vmwxUUwhycPQcGtfqMOt9273DcOuLRKN1inV69YvF6bFUxsz2ApJQP
KBAeONZLC2W8X2evfajOW+xRW3yHd6Rjv4SzNS8YZQUGsA2+/UwPc0AHtvXdE75RjlMvIwmF1YFf
mnaZjmW8hZ25eDFwVOdT0DpypDgM8dYDmEJYYu2aeU3lF3AjBJidJIbgY+lCX3c/BIwYcWzFqG9j
5u5Gm167pSCrd3SyQ0XlegpQNPL4jjpmptf/Hz9GwUPjUjOggcF9IlqxxQ8ZFFpCV5AXlUMHrwQh
lCLlZwBYCFhNr5Pk0KMImUyveSNCuQ29dmpZ0oF+56gUBu5m6sddUaBAqJic+5+lJ9yt9V4MrSTV
+/yij6L3V+bxToyBYn2fP3wu55B/6FDuIOwwRVT+k4Mc27t47AetQ9+2i2QFOyxUPJ/nOY0hEVRi
AZ+SnxxBnq8YcuOKnn9pt7Tw+Blk46Tc1eYOMa3qih19pemK1Fqpamud/cWPuLjmCCmyYwsmJ2yz
sskz7ND2fieYHMmVdwmaSQwEdifaEsjehdhT9AqUWokl5HeAEhxSVMYzQH0KJCnyKfYYjWMTi/jZ
FNlv87yFsqAmkAgfaMQTULocew5GPHA8OwZfQwTj4s0dD5+HD68jpEu/iSl8RME4TmNJJAYWpV42
O6nA32Mp+T307ZhwSuthhB2We2/8D0NOYYgBaccQ274IFN+AgM87SvrmWkk+2ZW29SC/CHIopdHX
0tg9DDPX2IwTbA/8O8cfwhA9akuvFlWKYQO5wB8q/a/dh+NR9S/P9qynGjapeNT6aPg9qaawJzzb
qdGx+h69hKVUaMh2qWoV6X9/UM0K8OVPdYFipd7lxPpAsSYVjJGBPtSG9kOTCnOClCN4M0h6lNPD
007yfudG1gkrVl7M6UEmy/t2VkQ8XlSxIrJoISASKnnDb06ldDDksRVi2oN71aoyVuBZ7MxGHV1+
k1NRifTRMxwAGFrtC7JiPRhVOMFVnGvGrFVHT3MA3eIHe+Y/wnoQfzwJKP/NxxY0ixP599prRbvA
MnByoSnEe7SSmeAo16i4wlXyZDFxj7IxNbolOp+nP0C90kiCZjXJK6p5spCieLFOAGBqOC8bPM9A
ABFJF1CsG8tnukpTiKkNKxKOAm9GjAGWJIpIsT/VtcyuF62ao8rEwURqJv/lQJxYY0Z6fV2KmboA
/As3HfZdPS2j/C0UC3hrXysFwZ8Zothu5kf8MPBeg7Ix06myDY4QRbLjSoSWKVQjVH9kBO17cuC5
Zjor9Hd8EcrWS/b1NQZY2IQg/W47wX1vD8qQI3Ea2yId9T9W4yjRRwSAJLyzkoPNjZ73x/Pp0JrQ
UrcPGuH9FQ+JAYC+/5ZDwkHpclqD49wyIyamxOLL0YpOaEIGmS31l74+CElH80y9xCeUCc6ChGyu
MZ8cGp3MN4LBKMR62dNirjJvM0tgI8j8+JLTsPmOBMetdYSrKLcOUrmYX68aJ4xbb0rHKtkLtOyE
OrhJhgBrBHyqssMapjAi4gjFu2df5vjQYiRtuDwgNHtfMPp1KjBvt7OwM0UOYp5n0VsXp0qe1awI
eqw/bDqtwJivHj+FRcHuApWPuHkF8EljSz6BuQ90XWoFk8TkyptZK57UKXG/cWmY0VapgRpTKS4B
k0Z/tkFHo31lPHMeQIUWN8slbis7SBaEofUTfEPxnDBFzMbNOm6z1H4K3txUGVff1cJe0NFXQckz
YiDgzzcjMDHLkZuaATW7ByjNU7TIj3Zj3jiFMciDKIUkhkvrZXM4p8xU+MmsSDuReIC32pmeI+Da
T2rQ9yP39PyBGHwSidIRGMhjo++1reuB705OxdWs/V9RmPzbXVY4/smQ2GdYtXulGnVR4Hvew4Nc
LvTCdlpNBkBKzzPzBfdSfIYxtbevFy18lPHMbvF/g/DCDfLC6Gtfb7LUIphRPFRHbJTun1xppy+m
icZ2sJBdDf2de8GX/Qu8FNy1hhByCibO7pP7xgglzwZkxHQQqo5pPNcPAhDgnGsBgBUkyZAq31dS
qd0As+1OHZjCA7nFqJ8ZqZJ/mvhnNzOOJxJzjIEvvHZjLQWEavwkAu9axUfdOHCMy97s73ItjKc4
Pw1jgr0jhKPye3bqzc/F5SYXJRyIF1+NOHyW/N2f87d5KxS+6amq7yU1dOK/TQY5rEDO35wuY4eS
nBFfY4JlXT6APet7uTSB5YJdOhY0R4ycO6Qm2q5IfaHoO8mRQGZgvpamKB1XpP3IPR7zwXi9dzdM
7B/gGVK2EOy8wRI2rpFXtD5zUb8uwefP56nceCXl/J0piWDom+Bf13QmlAOzvPOfHYhFOYh4Ns4W
IN+uQwOeX+DqDECioaFZ/h7m7XPTKEW7tdjicmv+RrEMMLMDBzTxudG0J2do+vu+fMOaEgoiMdJt
QBzLXtCp76HmUnZk/f6Uhu4RvuQuvWQPLjKSldNRo9D+NSavvxrpyvKgfbx/G/QFxYw+7GgktBQ1
hnxFF+0tdfcRQoWyMizM3eKSv0lTgdl58Pp4Fmcy8AOOD+H8kmWX2Q7ralXFVvJYMiXxSiuHa1Kl
2mAscUvz8njeWr+ZVBfCFlnxfiCm30r2oiZ7uZbbUH8fVD2kSUpMBPctUJK5cO5zC6bC4sITyGFR
JYie7J246t2RJyrFQoL+xf00mn4QBDF+jGcjRpaaqvMuvnRMc48HNaSPkgqWgX1WsgyzN+6wi8xe
rxZjKOYVxBXbREd3ZkeIRCp9eOd4Vi1r4tlKJMgSRYNZJxovbaXzx+iSuId813aZhP6JTWTorh5U
tUdjp0epdA6bXARoFsWyZc2FoUYgQFf6lX+EzJ8y2R0zTtKD61KOs+/9DpalBpJQhG+7HCmhEzyF
VzRXRz6rJor8z3OP+u08vhEMKMFNrX4IL/BnniQ2LEbRdQjhNKMhFeesKF9Z82jJ6QTm9g0B07K4
hvonJtKqNv+Ll7/UCnS3t0r28uszZ2F+iNaOGjLYLF+o7rQ6KsShE3wnR6G/mqUwQMrks79nALSA
h7a8Z7Z3x0Rl44gQPHjV7Qe6AryVANOLy6Asx1bEL0MoebjOH9pM8geid2MNHYcxQz/uRwfusHCM
EwdRxzd3GA1P4yRcoB+gQSlS+xZUYrHcga+9g4TiMU+BUZvr2322OvHUKvnFZSvMPgVyk2iLGYau
cFvvHm1TrXuJs0untOSdC1Vdi9Y3fgOvdqI2GodfLLsL1QIN0KDEOw6Cx5H4uF5ucxG0p6q6PTgw
+l3FZTmRyhi0+da5hYrlDCm9Jm86uGlRtQExME7KBRHSqsp/acbKtMLcTj3PdiL1xcrGSwrr4fEM
kIDrLjjL5HHrsHaUeCbP0YPYd3lntwlZmYkigtsbW+q0GOSjpmeUabsGDQ3ldgIV2w25EOa004Q/
IPy/1ypzl5oTV2JxRt0LY/F+qwjEbHqpdPgPr1yaDO92bvCWx/UoO9umaTqczcEP3wONZGvoulj6
X+SlfjQObnzBrmdxa1a53gBESYgC64VvQa87il2TnZXGNxg9gLkORjPi2lNVea5Sx1XmiWZWkvgP
LRAGxSNy995/NU8KSB17S7+4ZqCsM6BYfG1rezGbxkA11cGf7aJ34wW2dTz43cFJPpV0Rgo7cq+M
N543lcgsheuUhjLgOLf/OQN7LQrGuLo93XeCyvLAYZHuStS7ExlgBNe6Y/b3hp4h2n6jr9BW5Gf7
w5E1p7wsntPfXnho5zpKUXYZcyGL1rp8IshMTsHE5m5CBgy4Z06gQpHEy+ymDA4ENsFYupuRnn7K
HJY6CwdULUd691+ysGKHZZfWnClnO3PiQX/YbQibeWvr9gDGItM+RCGL3UpeaauB1KIImhg7u4Ir
gPrwl5r8cvh+hIMjfichC5LDAk0kwqKj/Vq7LzLsmelq9Yc684PhX+c2lXZedgN+E8gEIPKs8VNO
PoX2U/eA8ZrQiSC4GQ/GwxOxgY2enDrIkhuaE5NC/Z7+N+tI6oMpXbioqBNq2LQCR8Z8hXnYWQUW
1dkFo2tu/39dPgQez4DmucxKLz4T0dCmfrjbm+2bIKd66x9IndDkLRMco98HDLmuP+KXT8Zy4H3G
pqMj032UIsi4ywN/SArKE4KdvC3oiQ0kjIwj33qp765UUpxZZgFVzUxvSbVy0WXncUR94pKnXT6U
SUdjAVhdbpi1NQvx519pg3M+qzJBU2mHDezkKkjdVHE8nYapZDN8//VkWyUnt7NKtYbxcHwx3l9X
eDoBUZSc702Wcs/SaNFJP9ipS8Kxx9a4X6Tvmopt/maE1AoOF5dqDZIpnwKj7eJDwPhyJjN2K4ij
eC/CJXErY5i4fFwMpS81fZwD+knXT+cGo74snt8GCH3Ie/996K01IU7LanWijBL8EGnkZ5ZBntfY
s9z48uBgOVQA8yFa/vPWGLVdRTT+W8jTiRzAvKseZUqJxTXUpEtLqQKIlBsmgTMMXDUi8UOjPIoE
SkrpCqZP1mMyjEyXvwFj5YRX8rbhEGz2mK8Fnzk44cPyqJSPA5n2n/T0m7dyI6jVqP3jzbMYF0OL
+ITgUAd0LG80zpcMfGZ4XAY6zlcl0DG4TgNTC67BmKNNQhMIH6jGY2FBPI79Rbbjg585nfb/bsaJ
XaJppUy2fzQwQPHUV6bGNLUp0/Pm6Pc/TZxYcumSOMXVKJr1OqhImXoXYCf9NG5ce0LBgC2/fXpu
lRcihnnS8xKfLLIY5k+RmGO9G69LNT9RcmCNeUGVGngq7/a+4Ff+aBUugJgSVciyFN2Avkv8Z+6o
BpyMUP8YiR4JMOa0Husx34ktvf53my7cVRbOPEgILw/iQ5BTjhulG1wTN2P+opWs6WkT5S7i/aBo
RI/WkjE2ml5ii3pbbo+WMb3hGitQbY2ot6Q0zXrhEopEDqSMZ/DKDWBsTijfJ9Pxhmi+uPiIs7Ty
WES9vNbiK4RLaZwqf38jNcpbBeOsQ/b/he1vm/R9bHHrj1KkLzaDcL0ge6LIi/EV1n/Uq6XKa344
IHakUpX6ZbQK0d01voRQSdSGoLQOVut021rI1U1gHk/MgrRSi6Em4ihdK1z1FPfSpRmMrzdfEMXQ
ofI6+WQu5DxfxK0wi9WPv1g1cA3UT+3M4oFTxFd6Uo7qy3QwDDTEiN4qkkPxXlnR5FGhr6gP4rAV
01yW5OsKuKgzQhvwWZPbLeF15EQ0z3bMnQ3/2TjAdIaH2a2f2pJYKXVJbarbFas9MH16C3AyykQX
Qm4Tb8uoqQKVtRbv/dZyme3wQ0O4vjUAgJ6AOqwkGptnZ9nOSTT7Wvj2BP8bAAdSvZc0lsYBjRJk
GTIlzSuWEFtn+3Po90ZxXCjF4AV0Jff6Z5JTmEApEeLVNEvROF71cvexZRAXUMjjfbmlWxc//g30
sytm3nCsctHLG8POvB9ZrEjbP/BZ77NaRZaYYSLqHXfL1EKWHWKAvAxxAW+Q19kIqUBK/eNuiopv
2EIqvgZTnZbSSf2vj65b85oJ0CKnG6wBK4jsPjzkXeqo4W0tRoZZq7Epai6bw7/dTk+KQMHf9XKN
PmIudmB7ogG1iYK/b6KAQscMB6M8zIl91aHmugMhJAn1dJN8b9JL4DmXUREil1fHTx9jQ1Z2qM/u
FxodOCS0a8oXXDtCajNTCtEYVSfaYQ/mLvqsYb96E1ynRskNgxsTOegE3T8/oE/rOd8pFiGR05JS
8T+NV0vygdfs72FF1c/nF7nnL32VIFTKI1OW4hgzGEbjlX8Nc4DJs7nYZnt6+NzkEbsUew9WEAW9
Fil0TS76eaz/ziDPMxvo+aqTyGTZJDQuxr/F/RuNdlyEEj62PwZj09wxMr+4WzNdup2D6JvQpsCz
4YRm9Tyk1lkqCj9lVmVvxetVKiqxeLRS9gxwE3KjFKxrrOFSeL3MAfuaKu1z552v/cXwA3ESEmwP
Mrtr8wgBusHUVe/A9MGz5KjUkHx+sbbnsdMQncR89pXINwcjMBX+xYp/TPmOipRuzErA1JL3zYhO
S25MD+/gJsB48ZKlbSjn+URNcx2pTzz38gvedjlZP8tpuEp4rNjVLadhRuueU+2LR0GfD9Da6M5Q
7cVF7/CRGvzBOke1Zf36NFRnlvN9dRKAdPnEGjWF0DQwWZ3aMRIrHDWouo9rt5OVG9zDyTUoa5AK
cMpt7LjTd9ARkvFsX327sJ/Hb345lHOpBcA7v/xxaw3MbnX7chqWldHK47WUhe4AYaAwFFVH+fzU
Kwem8grvDShxU/WC3dzjrMB2JAGE6Z1qOB2rnQ4cwOfIj7a0wOsmUZgxQi0DTzLCAj8L1Z8A8Wy7
aJ3GBs55hPdpzc9YsO9Y9uJaBMEfNyvLckEZ5iiKZqC9RXUTowY8jbk3LnqRQZZPlWeO5QS/QJCb
GIYlK+kMBX7Cr/zU4fQnLi6t9B6aj55um3Z/ncELSU7qMMeyB3S0fW8AFjKo+6+KzZK/l9tQq7Gt
2Tut9ebPS7LBqnEkY4SzI9Nw+qnZjtkF5ihGmPqcaHqLVDTcOtWLi9fovppZ1KB8KVO+4zVMfFA8
QaO2omvzGdMmMHi/d4z1bzXukzfSWQ/42wfP04ZEFRGAgWCbUHNl4lrlbk1svUDnL99ME5qB+0H/
5HfFGOwW5h36tJbcZWQnEylnE28qs+FGpiEwE7OsY+tHTLlZoC8yOiV8qyOuGYohEQRDEuCEpc2L
DxqwkcYim1gZ9T/BUKQeDTvtQNrK1I4630TSd738NLa2W7nctxEv8qC4DsYDpvUrZW0h8PhKxLh0
uP4tvkHLbp74nyFqnxdWRQP+G/xO0VZoXOz9VcC6Ldt292ysIQMGh95dhQCOqOqxcZT+zVbl7agd
rA3cmt72/1tyqusDin41UpoE88cD/ZcIhf5/ud3vEr61p1ERB1hGeny40MnhZ1Babjpnbt4cgtZl
dmq7lbN3RG1VM3m5SiJJRKka7C529kUcoYOylQlYyPXdAK1aX2wtJRXv711iPIg0DWzXlDSx+c1U
uMgRWL8CAxRj9KZc92Hc68UBidh+2e/nQbMI4MAj6F/O11dU4vXvOw29c/VSAC9bTnpJU0fPHESO
NWJubdLTzbqMr933F5QDGCzA87D51fIphkd/uObvvpij+FS9S2KI6Rhm6TRQASIGworTTuxUrkHg
x0WLFytxxVJMdXDwIg5x4X3CjZfd/gBpeHnvnEMKj3ZDUCgEt7nxqK94SG/5uiMDh7Edo1Vz+KqZ
kpCYyhalQWpkkVqnVWPvTOIWS7hE3Nb1fnvlG/ghhqRSwQGT1ZCmyWvRta2hz2KbQlrV2X6zTXPB
jTtLjGehl3nBrPSFy6Ysd4YiwyYEwKIyt3o2nOs4Zy/OKcql4nuNm9wNAsvnPakJf7/xhGSIJ+5V
+Bhze586mwrVixpAiWvBTykoqxF4Ev3kYA/kRAV0CW673uuiRPsfz+ox4Bc4JkGK3XJH4MRVkEDT
ktFVjEVQYnLZAgm5dY6kZ7GOd97yLDiwwAK2pQ1RvPQodVsXBG79vbvfee+qTYT9mC98b/YX0Vku
tVQU/LJoBJ5hvZ4MmW3dcqpfaGwDBXlCM3JCe75jiE1SVhEVuY2Dp/9F5SRKqd2ecOw4cOjsVaDb
gEYh9y1Nkg+2sf/Nvjrj2yaKj+8mUCczYLaP5CQyf6LIMu8EGxGOqoC3U/Js/Iyyik/OTgoM3cuL
eZ0OQu3g9YrbwAitqOVQW+8Fk3ifzpBtNSOBZnCl3ZuF/ocQwHmVn4ZHIhclBiKK5U4vPno8GBVC
rRGM7f4Dy3oN63TDxGyJOjCTXz3qDz5gnDe8THosT6V5rM02FC9+l8n2+jWwZVoq7a/4NGwzebJe
iAeT9TwDNQ+ZphXOLywS4G8dXr/EEgZjiSXbV5jwbExLV9MCotxuZL11eTsk+o3sjxnRAbledHsi
GQc3fYVyZn0wXa36x0LrEkdpKPSLpys6qovqRrok+YTgiy3KvO/AkYF6cA+sgh7vc/mjy7fRerOV
EozunY9medCbVEFSb+mdDYQZd5Vh1aioxqzoMS6/d9ihTLS+LYBHqk4y5VlxxiLQnv1aF6cDHtWS
Fn8D8VpkIQOsD6gehV3zkzCK97CBuxERJSf7NFgiij4rgaBk9CGEQIfmZF+A9ZRxLX41NpqyzPRU
dT6Sw4ylxA/fn/2h+I6Zr5ePC7vB5e4zz2rMsLXLB6TaCgRJVwfVAzKkGerFw0GSpOAQy3Ro7fH/
DtwXjjEMBEdKfvJ6peh9smd+/RxQEJl4I/h11rv97qsdmwKO9cbvbJEJqAyoTQyTtG7xy4soFZu6
IRAWlHPXbdkDsYQx3HdoMlaRxxzJFwjiD8qYXQIHCqbTRmQgQLB6B1hathb+hMDkM++KUzMbyyFI
3LxQvRt1F8X9FUiY/rpVrXGWVQ/Zooe2sv7eiC61KFCRIYi8d7s5W0/O5quMqi621OkkhMwX62s6
ajXA27Jl1KRiGEFO7pz1tFMZN62MJClNnaEdG5SKJIv361NMvm9DpiPhetVcVHgQ9pcLTziVlWCG
On6SoXSi7WsVuC7/2xudci+goQ3+uMtNX80e2HY8BMOuWe+TYTuXul15BLXUVq8ET5EgRrsoiE7F
lIydPBbtD/tm7JdXFgQN0yamAliIGmMxIUDNFsJgNCaX7Yupj/2v9l+3CYseWazPCH9GZg3L4td1
euj/xoToKRvZdh1RiCPnSrnJ3RdeDT8YVYSOPzUdsKqCNFPxKOyNR8rSqtJJ3unwXB29iSPhV7P3
hZkgAoP97GQs8M4BWFSpR/vd5CVlD/e+KnIqCU5jah53l2wQba4+cPRRJ62ZbLOz28ybTAG22DkM
b+cxVn9LwRSTnkpyo6+1FPJ/o/aZy/amzGwYYAx2h0Xrbf18Qtp/u43upNJjl6jxfVFxYF4yD5n/
QDT+okLyEhdBd2LCEFzkvo8s1NsMSji7KNpKInnag9yPVN++OnJkha/EreVcVw5NxKeYF7ftb5B1
vwaFiJcXW85oUvUKmWAMDBar1uomGtnS4zW4FVnryURQZa2np7xXx5K4sRlj7Cso5Y2WzsybG5B7
h/ZcMJTf7AdCq6JCzzeu3N/bcwUdJdGleGv1MXBar3OHpnimhQbjy1VK2IBhgrvbBLUj4/T0BIy4
p9++iWOsJvjVGAAIGZlBurNkvjOCSdqOcS3xxCQzQrVgrNc5Zd4a6Ea0TPl6ST9FxeiY6eyu8Bbn
pRq/FgSy8H7EZMNdIL2ZL4//sjxTkIrMTVfTMrvGY5C130/lHyhRXk1QUDJf96xiBO+L+HLOu22N
fzIS+Ahn4/uiVwZekXdQMrivLTIUCDvzxGk7gY5Gk9IxqOx5EQ9/70GLbdX4Ou/51VIfCZHbY3/u
qE6geTff/zbaS6gs2ABkVx9Wk2+gbI3UoE/hRDdxdjxhbn0RvNG7TqkiL+uICf85slZWyMLyjw4B
dL2OcEosImQOT7nIs1Z5O/QhG3MAhG51ikVoHuV5fUK2wWfhrgv/Gt4nS+T6wBmxHmUAbxxx/jd7
5wm575Q4TeLsQmKITTCYHv7g2GL1jOJFnXzZ3ZsExq5Ad3KAlDPC8G11tALf5eYg6idITEZ+ToSH
Z2ucH1rar4sQf38arLWpCbIfxZ9qOkBu8sG8hto+TnfEhN4CPmRh7LfuiNd4Y2VaKB3cFGvMlHc4
0VQ0bUf2tmM8TYs59rziEqjUAvdwEgLk+3jUAA1NiN4/ngdUwEh8hwqY29KCzssDHnfE9SHU+BzT
rsUpYug+kRw9uBLlq3fT6u9IBqq3xSeilqujLpmwGLMQ+8aqbqnsacTfcyTXLoCEMZ3lBhBiYbLq
BRBT+jXi2ioxWeB9rZ5e5UaptxjyZ6KyaqhO5RlLMiZPup2EE0Qpy8GCKBtLhv+t0YnvOMC/MQBG
8Lw0gPxzmewSVxq7ewklp0WNpaZ4Y/b+ngLaGXMbzgNK/zZ/IyqAcE4mYC1FZebtE9nEI7xLGJOz
E1jRKxjSWFtY5ZyJrj2yG3uINVORF6Fgwm1lOM8whiklP5N1gB4ZK+lnRTWW5DRdvwIE5zYwLUv9
peKqIDMJ0C2PYHQ3WXlb4WZg+rYvLuUAQVu68gTB6TZ4Lek745duAFgrQ3ftl2ZghRhJg56phV6G
jn1ZmLSbLIVKEWg5P+hXGttS4S5ggu9V1eQ+boccXUbEu2snJ6kJ8aOx+RQ5xj5fR/JyyGYLiGXM
5d3sO0d2Fp+XFFZyvVtkJ0GoY9/WlEQ2+LQZkuQdw0BRaz8DT4fCn0+49DHA66Diur95AByH0GqD
UAs/eFB1WcowOrdqx2x6PmmZ+9mVSGlva95S8098eXVoV0nA+uzE5Snhf+SUgwii1Mm1iP2eao6p
wYSOjAOHtrUNVXL1Wh2xEteZir6UtIRGjXmtGvyaZGdnJFxXy/ODruP8OQJddo/0XKJ/E/DpFvLR
yLdbimTpUvW2/jw0PsYHJ/DG2R4mXLZu97N5aSL2RLmeMkujx33P0H69RJngFWRqfFmZdME0Y2MB
1XlKusFf7MqwnvCky4Ny37uC+x3j9IYifxI+1d8k74sZvRMW/LV0zqdLHtzGUz7aU8UHw8VnRtsv
NyIbcIp4LAFb4tguaXQkv30LBcSudrYMOo7YEDifbCWqWaiG0dt2YJtsxhKxW2giIu3c/ezmQqHh
WlMd1whz5fHTrCPNW9LletL8oAj20ILw9tN9mrSwDFqFz/LPFgVwbzAaypWvLD9uNkfTIwwLZJsU
OcgeLzRqtz2mlnh7RJfivV5LBseNKA5vmB3Qpf+TlKxL2LMB9sy0GF3UzEEstcYpOu3B7IB877Ov
XmWy/LchKB7wuCFQe8/pZNBNhDfRkphCWfp94UInaKSqvL0ZAz2td30BFSG+O60s7mlxF7lgXhAl
Ib3/ruTuJM3m4uKCVv1pImcTbOJyjGQZr+caBtAk1x1Jn4tuQLmgxGwYVnGZdgKBGJoycvtCxumh
CkwBthTfNlvgHviXneO1sA+eWja83Zra+Xh06qaFNbokMcR0YFUgQ+XGpv6dYnsjbOEexmwcVEhg
oby8OBla2jl6Qoyp2tO+cpwhV5Wsh1vJ+aKVKlyh1fJVSy/Fr2naYmJmlnE9moCJg5Sfo23KIZZr
y1NmI/HIIuznbFRiswXzVRgTIl2z9qiCSLstqmMajUjVOKL6vQ0y4vGLofDOFJK4jhY0sNr1S2AE
VjsnEWgZvPNp6kzXhqb4wWMrZwpqHn5cR/s0oIYxpXH/5JL/DYt0Y5OxD8mKZCqNNr+CP1RvAzqE
cKlL21T0QH6AajRhrHQdprJVTv0OG1qqpI5nKqKFHqvbm6+2YcM7u6fvW8ETSIFQa1S6qb3qJMJU
x8CxSuySF6pEwYuFUrPW5ftUkrcRtfT8aWHirKSSRLab5RD/KJ/pwrJX+9/vDHSHmgzsES1vGpRw
DtkfQWgmtPwTJYhbHkJ+4u3NzPnDCJricEncOXIzK8i49m4/NEMkDHx5wlPVHsy3UlT6UM+79jvq
t3zVuL2uCIL1JRwuDgro0Xay1GQF5OTUNcBOFHWC56ptPCVxd/9yvsuL3X0XWJarnwpTFuziFWk9
ezzBGNCZ5f7Az3xxSIg6cplhjsYfaubPUTY9BxyKVpOfaOIg7SrlJS+pTyOfs+9hdwBOSXT6hbGx
DXp+fDjIuvXy/OdsqVEh0+5ic+za0iQXjeB6h30URQt2R2U/uF/PyIymFF6p3BveHe/Yp1lK5zoG
tYtD/5dFafZaobCu5b0wgyZ8BDDwq0omkREZJWr2U7cQAOxZp78KXd/divbhDrjPnHbDb2oP/c2B
Seus27SbqfYxO9fqJ/u4208MRUk5W16SYCTzlQHRzUzSS/wNjjooEMsyZyV7SH24xqw1CqsivdGf
dnb3LdLEE5Rvav6ZJmwmkr58gWyG3I5DHC4KLORBlbG916Sx7SYDfLdF7ISUdmh7Dv7tnRdp98gL
YmPOo7gZ8XWOwZKmvkhW8rpMUvSiC51z0qJyGnUvgwFZ5Ya5XKeweT5zy5KvFwy2VFPB6D7/wbJq
a6c7EgJJ2bCCmQ49sO6DkJ8mIwgfS1JFu151bk42zsslTPTKiwRrs1A9ldJ+5oJrUhOaYZfxR6Gn
4ixcGHQpmiovqBOOxGuVI9YZQH/Tdn4uPoo/znaLoqRWVX6y+tzhujynNGgf/5b8G+DFdlEikU9X
w+Gp75bZuZZsYjhPlfbsxk+sQsDKZvDZEl2PDmmlFc9SIGWW5m2vBNq1zOqFD7QTYC5tG1Ykkv8X
4AYbgElMehnFWJABkLPbPs2aU4hJYYSwSc0s5QYSlhs/mLlIPAujV2KPlBpLg2TnmrTtYim8/m+D
hK8q8F8JSMaE/fcqzttSPIhdNThgBp/U0n4nkjggcrhWINmWwBn9puLmla9Ei/UR4CCG0zpIZ4Ou
5ecMZkJIkbYAEt2PuCCMDs7YJoMEbRYGah8gVFT+XW5ymSS6o9lIKkKfwThXL7IJhDr5r1Q2Qrn7
FIenMBOg6QNuoDKBRVdzoGApMALD1e8DnsXZGIsLuav+cMRas8vf8uQxNRt9KLix9waxajmo1yka
Kj8JTGrjwE15EIZ6ltH9VuZbd3t4uOZ5Ocdk5RiynyHFaK9K8wgHNz3ZgWo0vdrgUV3D0aGQj1Fk
ybdyt5y+Y6qEy8wd/0P2mUeOGC8+e1P9Id+KqIYeGmgZLxUYWRAGTZW7yaEV/Bj96ves3k9DnvAC
Mzd6GwxkmwMSrfvtK7A4c6QfVCijFiLIQE1xeq8JMHOneUHLHcCDrq4p0SYwFOEx7N5YYGnV2MEG
r9+pCPq12IKSR9aTMHpnp6w08NMMSDOOT7v9rwoUms4VxhWL37kHlgBuVeplgCnN7vPLJHoSU4GS
XlGmPNf1Pjmkv413sKqZ6nUGMOoKlwUObWfb3qI9SqjKBWOQQl3HQnlea14furjHox5dPcM6Wn8S
3FlFVUUA9uDTdHk2i1c9cLEYgQk1FMWFIEEHJ08qoJtJ4UbKMK8Ed1dJwsoz9rL9ZkeDL5Z6YDrm
lceSruMdRrHPFLznCxeV+GQ+n3WkY/+R+gtvGSiGrLEiHG/fU7CZM/x1BzRGZPZ657s0Bzv4Z1ep
NTOfEilbjjlaustOiFeNyfi5YWz/6lnuJnhTdPoPZ/jzTzbTvMQSuq6P0I9g4i5XWiucAqLv/bGx
s4IWy1HYqTu2DwIPnJ9kxEGpnrUjj3zjMbmSrp/fEcC5wNInBmE66s1FsV3p4moFfkhFh6vjAUq4
CizzfxPv6fca9U5DnQdGQOdzJux/pn/AaaJOGnUSaS1Vf8K8GwbtSex/gXsfFuWER0Rd86sKmGbK
gYC2IGye7aEYYFxnGRIP4tQ/y5pwX7Fpvhbkxm+rU1uaRJXCS2rIK3mCnVhZGZfT4PXfAa7YJmxZ
4UQnBMhfNwMdatvwQy0tZZxumdY7aEJGFtnp1P8Z2BR0HVg+EXlzSRK5zXwQl0S8jjGzq8bnnmRJ
5IETjzwT+LZEPtt0VDkZukrnTJ2kvNqyh7hfK597FIb5KXIO1wryhvJNi/778RjThNkcvnPBZ9H7
2HzWiqe+P8WJAg1ia6AEU/VDFm2R3KtAkvG6cWROaWKtoNVlUCWXaEbFrOv9WbAlM5hFeoEEsRdj
dsFjG+gGd1OFcMqyOaaTWsRTCBSdCmpJ47B+YV2BaRSfgVbmXPP6aeAb0YBsun4BO1oWbWTGtgnI
j0JGj4ygJcaM+zyLhyYez2kVblPx1pP6i8VSuApBxqHQKQfLDlhtM7I6Nl5/u7GwWeUOZ5zKpWFr
jgSRz+jtFC7RXLpXi9FGocK4aZMw16OU8CdwPlK1qZ9JvZJKmD0VmIkZqWxi5NvOti6AFKFk+qe3
90cDZ24vI0t8YzOvuN6N5+3mHkAKgQDSD9eG2FMtSw8GmK+Ui2Worc9nmYe/Kai+6c5pDeGDY3io
g8tSVQN/IZXLVciV8IeUmbRQVAsQZTtmus5RvFVr4zWuAMWl1jKvAckJ8vDZL+61lvfNRQQqMjZp
c7Dv3bptvT8ExlykZb/VYSjkP4d9+MWgn/gbc+pI1ysquXfVOz/MpwnLIpInPcoKmZsXhnJAbxqo
qHt6qLfR1PqTXLt/5WlfxSMZteVTFNMT4JxJdC0EPvJqKO4Da0e43imOiDdVMyM77MqTJixSS29R
/XFr0uK3f3s8WHDfx+71NNBLhPbfq3XwWbR574obq6Q+MRNRRsT3rtS8uil2I67vHgHnwa19Nn8J
mFfdbxRmbCU5nTibRuBUN9nuH4rplCNW5L1p82r6Er+UO0XPjzumiMvmuMWh025pT6OcBs5RvLdU
GhN30h4bUVEtrEsXvM4WgmkrW+5q4p0DuQWMHLv6AT4skOCIllXS8xh25M2bi7VwyOiSqCBuIWfI
YzvCv8t5+gxpcsVDGfq7OsetFa6XVyGirG0xStAWUzqUMfdEWPO4BUxgBBDiIO9RtzVZ82CWJU+X
Kuz1Bkq6FozNI6XECF7Ucnzmy2bXuKqoVVYyGrZ6xZwi3dlfYNTIi62dgLjdwrPGzyK0awgYtO26
b24X4Mn2LzsH0G8Qs3G3IPLtDYjDa11zMHWcUagk0le1dfgJAP4VQ7d3xwQYWym9zK76WJlRc1h0
A3zvamVTyrrso4lomVT8zu2lMR+IFF3WdO81CHXltYDp8HYm45CcmS3B9zd0LNa5o5Gjxa3op7Vm
tUOXQugjXk4dd/LcKGf+UZOfddhHeeNRJjqRocQE/RJ+0jQ40zqB5PVydssbccKtU2M3Pv9YefuF
2LG8Fdw7e04BjxtIE4vvBBrItyzQgRRzwvU7s++ZXvMwgtQziS5ap3d2L9AyHCxGjkHahWM+Gttq
WLVIuyyCVv+eyFmztisVXQ3y4gWASCQyCkmbDIBAq0aMD/TU9iPQrWtMCZIa3wPyzn3S5hUgRkf+
1CtOVctGyGkQM+C41plXdBjJmDIH51gl05WcaXnnzIExwS8aDDWy3+HZYDCA8uvivmPeUVGV6Fkg
fCCMchY1UejWPfrxrCknHcLaRGaSKcjDHN0FZTxN5K+s56O2ZaJeHAXK0sKEP/2hQC32qk4Qkv7y
X56gqAkcck3y2wwAynfnvnPmyEJyKKLWYr7Br+hmJWwB21agpaLCgxrJyZ9uMvs4ediaCcFO/RgT
QSKAJCHKHfmgJo1KXFXTlk0Fd4QogJyWHrNU88W82P6IXXe7g9LEmmrRdho3TuiEfh29Kl8G/VvU
sKA0OKB8tTSTOxikiDdvmGynKmGMOJ/4lX9orru7O0oEkbcoAVEW7saraqyAoRAzY/yA6ykzoO/o
oXrFIjp9rlVV+fZ+1RGVUlpVIN19b1n5/iHfPE1oHXD+vphRY8ZgFnPdgMdS5R60g++k4CJCLXaL
ZfOtAmUN+0hURfstn3quu9hySnoYpYcxO4pHSHQVvb8yzuOFVTAJuMNuMkf0UyDxigE/8HCbiho3
I3O4HKhg5OL26I8G9wM2C9wJKU2KANDBlmUuOet4A/7YTmeFLDAobPQP5FD3NVPWXRf6HkhgTC9D
72gq76/iXYqDMepszLTjN10YmzvawP+tSAS2vdQ+2FKij8zlZJP6GWmsg90RZWay1Un4I9OWVnLO
PTLlww237FiXK/HX7ZcIwnnz4+fTHbxVOaxiKPMKHorBkaYqXzxJSZLmuHC/JD8WSyAxffpVv1NI
lMWcc5CbqWirSJOpYmOD2Kzxr5LVCcDq4XyZOMR8ha1gswzrc1cAajjmLkvdoqQLaZdnOllg9hIV
Mw5mGJpTc7CumEtUhq61Nm79k1gmbljdmWk8Ejtb6iUwjKBV77+z5L8a79fBvsIULsdN5z9Y5ZVE
PRnOsGYc/nGPkKw36spM+D8EqX9n0AH3+Hv4NJk9spmsRe2LtRtT9FX7JJWrzddRIjopfop6EhGV
nVSXJ7ebOj8jOF87k+cUVGyUYqehi3tNpKnjFa9IKubMoeDEXi8TJmOqNGr0L7RghvQ7Cjb6uBCD
+0q0oG36UET9RcAYNfJGUfkHxGvxRJJLS0201PGbS+MDG3XLQjdJ68H9+NZECeceWUbi0APD+wch
s5PHpQS/UdtaPQ3UwKxUDU4hWhT59DqPk9XaBqIvfSyqIqg0yWE1pcwuZYnWsss7jviaurKUz1sN
wLq/P4AQdzA5ktvPepcf/YX56cCQGTgQ1aavVNzNmPMoxnSGqXDywA14TJY+7lPFUfuhzWnNct/x
JK4f3ZjZOF8fqSly6DwP6TdkZupilWPGb9AeqX57sSMTvb/O1nGVtwLr8rZCB1bgKnF9Nljqa/l9
I3ALds19ip6ZHBovkKWnLi4lQ+en1Q/wSgoyhogCrfiaqMTuZCxryQVGh4ipQp/wGba9VCII3sjG
hpeqx+SwpBG9nTNA9Zy+G/0xJh5rKS+KLe+Hx/2+Z7vfJI87EOi6E3Jf9Cll6oqQ15CuKQlVOMqj
lIKDLGADyJ9pF4hbGiDQi20qeROfHdvA3aITA0AckxQbTco3Bo2vlTQxThaKtsj0KCshtYjbRU4g
HQpPOZ6Q8o8eJmNBA3T37tXsIb2SOhd+OjBYZ83+Kmqy36GmAhzhGCAnUduL7PF2U+nDgLhTwveb
fpXPz9eFSF4URzylM0ALC3Lc3ZMUe8XP0MHJNtpc0MIyhJccqpZP1tCV1hAIb+qVBUr1Et4CuYka
trmFdp8QRzx8QdXdFJYcefAOIAyEwnIO/uXkzsfCyIeFNNeAlRamB579dU2cb6s+KjQR29lHr8e8
VmlUUuFHy5vBOyJSEO8cSOam1+IrpcM7aPLq5LKuqJzNGEOkhq4JF6pzPY5g1oqIxeQPYiFGlWWn
V+szeOo/7DW8P+iXD8tffbx+mV7T58ZgILr5s77O5VnDDT29KbTc5eVusOCz0a+DEW91221Yn74Q
TAT65NHSF75/yEo/lEq5/uz3ojQGePSZmTYZ60MP7fd6jIlif+C7Mo5h4Zeof8u/b44RZ9Zf7A2D
c7uTCVkpSY575eDjYtNtIF7Hfech30E4nZ7pGFxnoZaKd5EcLykCy8KYSVi/RGdfAOKujPCGvpCw
Xr7d71zco5z0v35CrqykalRDACA40nTWmuzB2kK2+CcfPwD+C58R5T4FxzQBsGUKcZ4DrDaALXd5
aOIFx+4Na0ulvtOOaJPvwjqkyWBi7T0P/KRUNTy398FPqnyjvzdfUxTIJXZB8IezCZ0bHJHCOWid
XONlS/weQZSDE2dGplYrfoIAuB3XO7TM0L5CJesxy1Ybubn2+iK31V0/GDD8J5emepEuv7JgPuY3
jphTCM7ol5QqzHMXYCzlhoYEqGvGz5e5Z5O+dOQl5y485y47pV2R3+TQiX/pyGyFhUJJ+5RTgjEZ
Foyp8cxHrQokAADtdR9/OknRsT7BYvhK+GW2eAkYE/BtVyyGGsuzAtEbHOPlXE4ymDU+1a+Rm2Dz
g62RVLTBz13Cr18jfZXtT9KvGr8NwockW3cXNklJUozlEE/vJZ74wUAJaJCd9AVDtSuu3Bupg/mB
kGqMuAJa4ndO7rGE+Gwha74JWW//q5xhsRZxdHQVCnv3RkPeWQP/eR6p1/WNlanpiT+wPjEzjat7
TSrfsU9NNu07n3KM6FPhjggtbHYXuf4EGdsQmRWyVzCeMO0HLA4kGXU1f6RuvYgsy5fbYFOD7a8f
yUhUtn2KePYBSYF8tEznkoSHfUKN+XHsZtiUBlUv7kL4OKB1aq9iMfLW/lqU91m+q02pugbHZEx2
PNMaAzWP6PCVcAzRvv4HnuDkcbRoUNP2HyKcxZPr8AUG2WKvmhdcmLxwCaanohG2szobTZQpcJFd
AIm8YYEsutPBIX4icIXU2Vdi8rgtO2/ZpLSdIfaize7uEU7vrtpgSCgbrjBl3k8mBFqnmwGCmz8H
TA02/GBYVpJfF82K7KhA5y1fJqgLhzoiI9PFTBtSZ8zV9ECt5wc+Ob3Ys5lGQqW9/VcIJVNRxqtB
vezjAZu6Y/o1hTRuEVVj+IDjF5X7x9ebW0RjblR4jZifzdYUyY+EEBm6bFJ1/6vfAyJFJGUHhqJd
VXq/LJ/ibnWarExzR28O21OPpKQ7ZUK560sTX9dJ1a4m9/s1RCXv8n3ZdfU84UVWProPAlokRlDb
ZLnpnr45Jh9ujQdxWrms7o6cL4wL5wP3tyLO8xeQuV9FoS5PgQIxpPRQOJ6te9dcjR4KplN4WhZv
w3OwVtqjuHhxV4k/4aZu6Mv2jDE/a+yfbIzn97AKWv1dvrT3YeRyclGQXm3nLIzk22n3Re3x2gVC
UOJSeZbtJtkqbhUtWNgkAzGNLvb50NmrqQdf6bVZ2iI7tnT0fzactawmywWbZh6MAaiLU9NzIdZt
PPGkWekIAqaQeRUsrdc72juQ4/fF9fPVZf6PTJywnNs2VFrK9y5m8yLQ2saL8F+w9B/n9UuQXzp+
WLs/oT4FLMsc9SkfLnPVWKs4MAR2RHkSW+R0QWkE5z8gke0f2Fp6wcRS5mm8C8mS7HSjG/jEkFiq
p2yhUEBl23Oz2xmZLxqNjAg4ppmZUQjFwX/wKk162nvHatIGqSvAH8vEdG/f0IldsGgGdSiCczeO
+vYD5o/sFJomi2IP/7wRznM2vpz98B0do9SNDrs2tfsjl+SrErIhZ9OPE81FR/fdY2y0zzE1GE86
zyC2FMF3BtoyIN4hqSaSJMHLr8wvNdddsoZiRq2iCVpLc1bQVIOTgTHN0edzLfp7bf6GHFi5n6Tf
fcCdvx+ZxH47x+HCaebH1we4VeX6JTx9OBFiO0eE4Xd/f87ZKRh6PKueeXq8epptyIps8BTMahAt
DfxlQ5qIEqazF4jyB5t7vPyShrRjClIy6mxCztrknqXwxU730x3ag9KtiPuUnKxYLBPUwolcoNkE
DKc2pQsjMFYjVOisG52sLjeYzyxNbY5Y6g2BRKOm7JBiPJDCMs+ZrCLCuOwO2pFFibC7/1Jm9/tU
KtYIW6xHzOVgA7RX7nu083sdaPkkg15k1Bn6NnBoCZ3j8XhgvfbIc4dUX1f8TUli0o9OCSSOC2wY
h4qKPPp+2LFF5wn3sqG117SFgJu3afElFndhxvp48gDMmHoQiVdGapFR08pD4zVoHmEyYXWumGvQ
xK/9uzvIYE/O8u2rR4TONbuFxrn4i62k1DdHt6jl1iz9f1rTBX6Qrszj1wP8mJrbCncu/tkLsEYP
Sx+aczhF5n96MMEWHeKV7Rp9pAiYukG2swkjFjUAK3D6fwakj0dV58M1ZxC3P+ftgI2AIGZaU2Pv
med0Sn0y+GVmHAheAAlMSWe9XUBujktWVaqfxWZolKuZmh4HcuUSaQwj4jDa3IvYj/rKWBwyU2bv
nr0IYNhJvUUPZEb3QGZl/PO/DVZX5E94m/lMopNBcaLcRhmFQFcF/fiZV7MQDlmz+pjN4oGIYp9d
ox/cxfk+SuTs3mD+8yeQLgI0OCFJp0HEo1gkPhuQIsOM8SHq8qyRw+e7r5a/j17hIMq+jBisps4U
4oPC7Qb7CXnV+YyLkcvMvG/I54bDwoj5OspCog2k5argucR6MzfCjDVmUCv6tAOZY6Q0TRWDyxug
I24gvnDYmL+p5Yto9sFZK6WBB8qJza7o7ZVyvvP9atRkp2WRcTZyfcN0m0x1WWz5YB+sGwbwDMT1
WR/63S0XvFdAQkrJCthTWuq2g0wrN+4iwPDy+8Mx3W8PGhocQT0zXLsTkhlpJzSZefYULRcP1/OG
GZt+kLTwnXk7/XUkhbNfTNRwaBVmoxX671NOcmvbjTp+H4THtxkAjFPgBKT1zlh0E9VzmxP9Flcz
GOM3YLJChs1/FQvgsz+u5lMIZgxRuWBmJYrZzfTk2MVK1s4ZONHeDsU1xyPgZT+hiV68x/P2kmXg
MlNyGLYVsyZk7v7qGaWLpjV0sGHy51xWlFb96Yox4UqLc2XkC3B1uYsgbpFDYaZTk/ILcK2t2ba5
oHvtjvVs24SxGnVjniUeX7oedBdOx+jnPVOWnjCgHs/YLQQpfdgJYam6ke9gbIT1EUUz+36Bc5bp
BFcJ7+btCkQc9m+Cpj/ig2E+EGeivUT1rjWh45VwscK4nWqqiRFs2CU0vBRBcizgPzDoRqTI33rk
UcdklbosWiw85UG5Hc+MzrRJqSf+s5d6QVr086tQU319XHEVualasbmd9E+D7m8ulabi38DxCSY6
p8QUIzjf1a7lwPWBpUxtoCEg7kn+qswbebFz2JYbnnVb/mb8wX6W0YuthutWhSA+uKIaADinoh1W
Tl0oKGYbpPvuwSxfhtFzXRtMSXjalzzdDEb/9M1dAovc/2g9OfEp8CeV97TJVI23D6CRW2i81krC
AdR/1foOJZCpKkrorPpXzvC+a4c45842tmPrqV3M4bW1ihUOuu67f7x8Eo9GcCV4KNSBjhvRivU9
bFhZa9ZHsToC/oW4rHBVRiTqpQ8FXL6G96d0Qis/veHyvbKebCaC7TjHULMu6o1O08rB136tSYUI
ERwNiQ0H7ZG3IaoSYh4NW/UY2Gop2/dIc80C4LfqDbEP9QltDHzKB1TN7VZOQSn2v4UzmwvhNKSr
JxEMk+RSpq4IvJqPIbXy+ongbdyNSOtI6DpT+U4i1rmPdFbxXYnNJqZhs/f8sZhhNzhDQGbmwuPZ
9vooHV1+dNnURyf3xjdSWvOzPH3P7FCq5j/UmxUAHnp4+7J1p2mCZNDeNzx1IeMiDpqyVIKIevNU
FLmrl8LdwXa9ir2la9qgydGF5m7SqLn2L3qgGNIwKKdotgkl4h4/8Q35Jeq0VDOPwFcciNzkz2RX
ryR9JHCV6SnImXAzlKVamyXVv4Am/MturHlmuOmfJ+XvVoLYkB613xYS6pN3PgUgzjzDuaXnfdKP
fF77Xe7AM59KBoLO+H6hGIhsL4fxM8+EKTwBtdE0FBlexEdKU8HIpbpC/oLdO9UXqFCTAQ71M7+p
R9rlvxMM+YdwadZWCBgeht3OsenA91CoZdEmis19xqfERSLbY8Sti9sf8Iv0ZLKLPnI5lnMxRYus
nqiobtlvu1aPWuoZ5T3U/PtuFoJzWOmMPIZOd7dZ2mxkanMnxblfSFqFgJndthzAg58sf06ZOUgs
dxNRsYIZJCsFgEyNH6ItIXo5Ule2xjS6R/nMHykU9FnEDvXeW5ptP7HVcUY2I319orSB7XUWJAd7
CVoMniU+BWx0SDiCrwR6NhDBiAkABLmf5VtQCJhVgSm35IMCOC52OgNJQm8WQEUob1PvLXu1QXNW
3uZafbw1l5FAC8+vAdOqmS/MzGJNtIXR5V9cGwI27a3gDx31yy8R25TWevoSOL1dY+NBgcZHQg/Z
njNIai++NRH1GfJOZeilPb79EKE/KQiScvLg0xlwULi4icQfw6+Pt49F0jznQ4NVHpEZgyNylOTi
0Tz7Dj8PXG0p2yIUY4TV3F13k+McTxhz7TjzU61b+x2cpmjnZZd3uj0ABPILE3oP8c3QT5ysMrDz
qcf1DeYIvgH33CV2kgrCdpugELcLDPdY7B1ar73Euqa28f2eOIe5/ONYCgcNhQ+vgqw39Q9z/tF8
x1KNpPYtyCx3UMsPJluGooQkuczLqnsJoLgAHtyjH6CyOxElrrGeVvwU4KhJonqdNDaElZ4aqVn1
NoBZ2qoOgpsCV+vcEa8IH3nhc5iJxH7ucAwDoVAVZRoOaBVU90+TxdaxGWOSXm5eKyuHF0bybeKk
CvtQfbzEuIn767nnU9zU6Avxgeg1aJfX8uwjX/GYJh+rsmubkVlruiPhOqZh/OtJWxwWFdNAf98E
kxnuRlVqb+LFDYmOvZ1aWYNXV37bob+z1iqs0/dmJ/flexmCcPB3X0YyPXpej0BE4kpzyiEwFNYI
XwGAWO3+B2P+m1Mr1FaoymRKctFwAqr0iK4aiTi3WmzqCuSW6JIEdmhKIpH1sWEuLzuZqgGaa6xQ
AEbu/GMMk1IQQI5kubZt9PbyX2awRK7pSWGnlkFanD/4IQDk9+Mc3IqTm24qnfnUH2l2PDjFOcvR
emfsqiLxsskJzIKSh7MfhkXQ3GcRubHr+nODOruCjZUBR3wzUQqkjHdR9WUPSh9YCipSi9WcOZeT
0AOp3CRqSMEDX0q7+mBiuyTOfFEl7JaDAnE9U+oDL+zMDKxnVViBTBi2sasID/rBwSRRZpR0TJCV
2wdOxRxbXM/L792cQDLYDdXwhYlmVNRSCwfrz/EPzBeXoB5rncXSDHVr3QFw8cwMaL5X9921alM1
a1/+hDFbLCERcN41JvEedvttocNdP4MScRocVJHEr8xVSNnoNXJXX9DyT2vGu8k+dYWpt3Q3sSmB
O4nI3mhHoxWUGOq0XZypHfvlZcxetGrOGAn3huLRyfwGJrMS/xdd8fDg8EN7m6PJIPBI5ZN1KQtY
/rRQsUlvz8BWoIhvg6+PtpZL+GstcMHaF80Dcdw+SoI0667OepSYu542HcevE5eEkRJfzsX0WUkN
fcdpEDifEUkHGapc36ZGDxgl0ksnplcIo6N1SsYiVWCrSd1mDWlddhdEE2rQDr5PhYELWKNL+tvB
fkmVyq63wth2+UAFPIHubZ2kXFdDPCQbsy9ySvAvXfSPfuILjhJ8if1VHbT/eQy1kOCNkjKb9uxj
ucv0JsxvrTnQZtgFulGYs55B395SosxOJGeAv1uc71dpswINRsjbwuXzzaMkm2zgKLrkcYQzSNpP
OXJww7sss0NH0HcbLDp3H3iqo7ywq1bQOjW3vNkleTS+5Lisdqnvt518kuiogRExwWKnTjCx6t6v
lv9ARWOAgym9mqweAPe61OAvb78lbO8d/bAf7sDa333AYd+2ce0kscVXeSbQGsV1RJMHhdZLErGz
s2Mw1NVdzrW1/fiAykQYvuzlag5+wCLdzZpEmdRE4mPl344Q4FSFEEAwrdiTUBuNKtfnvFud6ohM
3JITj+wSej3WviBXzKFMYnvj1uR5VF6M7BOOPlUWR6mXpf+US8BvvI0n3N8h/UQjPB3bTjwHV3Mj
ptdaN6UxMKg5bPq1OmfQcYmuCkTXd/ssl8+M3nn576wkcxJ4+Q5rycFEd+19mh910+/iLniU8cpr
8vSTk3a7fmBx3jr8T4v0+fr2FenAZdQDx/eqWWsbeZ7mN1BWqFk1WPd2fSyKsvj9qmD/cFAlPa7L
kcBHP+eAs1OgKzVlrpvNwRZabVupteqeiCfP46IspkWXBMXySK79S3mMcP7g1YaHBwCNNsR6kCha
8WzypME7Tj0X9zM1aE1JXM4FzRCrZZv+yLTdpkN63KPlD83TX+xJfewi+by/f+/2j425osWOrMjg
NU5RcS5MzU11r4Yikt8VbMV0Nylib9Dp5POrANz0MzyWh47TB8VwQSIYHyt2GCYG7JX0RVTDl72V
QzkOS91lUVYx424ZS0v4677XK9uZeIApH0cMS+SesrooLPOA9XtkIsqJQyHEk+fUfFGUsSHyOxPe
DF01gLORiEICf7PEwY0+XanyFGEQS33GKi/UtuSjEF7sUV+Q/wTAMR9LHLoxOxxHwHfRb91jKb0Z
8zGYw+Z8QtiQouuQpeHnPccE1PbqJkq0DLA/w2Lgs5NZV5wNSEsdi7UUFAGU3HNXEY1UtyJXK6An
9uMOm+eSHF9KsTLgTeuuEAlXCr7+rKe3SNLuER5TdE3fybofJwc7rp+VJ3XUPFK62esL7Fxb5Rbt
tKOBBe+A4TuWevMGMBnZq3fv1c6c7qzTgEoMIImEYVs1fPKTx9yYkX7mD/PK2YXzCgGwhLPOFutT
CdSsG34/6bAOG5iNInXRsT8lC1qcA1gY9pH3ymVoHHzj24afQBUYAXAgkNVWw6kziHuCZ0UacXbT
NsVPDHIIo5z/9xTB5J/4uigOypnIZwfuQlS3jdLDqO6cVVZmy7Q/M14dD5gtPhBcw6+hQjyE43QL
6dTrXtt5di32WqtbA6gYfjTwFalXvc2lLHeRfjig2veVmME5XLYWZYoYAafRTbiu0asfIWZ+hCMz
h06GMinHV3ErZ9IUrNP1dOVoSBpi7rEVgBpUM6MKDSHSOzmMivlOTkNQC7PNQN8q5YOeKFkxYuPE
YmrOczu5mJfP9G+cWsFBPiqFOI06ayLFGCWcbPxe+5aKO0GKHB44dOkKatRqsJnutQbXu9rPKRyn
BlbtPiF8nCZ6In8Wva8JdwimI8Q9P+/tS11vlCpPe04wR4hVR/5zFPKBxEKhyGe2QjwnvJ/nC5yo
ct0yyrSQo3bqUl1yD21QmilVYRQWBaVdgNxzOuaJYUa+JoQSQRwPNC/q2odUKytrw2XrbiU2GxEG
bpTaLP/1r43ZgBzL/RiC0nL6YBtS+D1qmrtHK806suyWR0/YLa7ODYmafoDZYzNH7Khw7NNKXMFF
nJQmX5yaWl0O6o96+PGtQ9nRbX72w+wIeqC5HYj3L3XdBvlv2zloDwpdHbmKm/+Z4+fZXwCtVWTF
IfFwYIVCDzS7TqsmBcQPRyHwEMVM0g21z5+NiUpZj4nGLZJUAsSO2LwxhE6DyFDdC7IW+Okf9OpS
CufO2iCy6YcsHNGufbH1szikrlD96QcIbS9v4WkdeTzggm/L3YI7uAguqjLX3dKSlA0f0yjlJDC6
92q7D8ZXR758DcfRB8eOueh1EXclm1ifvy5xdHdCQVD8oc4AsmH0D/DeHdLVWGNC2r8/exef1TZk
/HWBtVyYpH2XJrM1mZDzKqSCrwcgnJ8N7M2332dB8aff2BbiycJ6du0spFAc6FYAVOOa3G6Da3yl
86dHp+Ustg0gJLbJBavnNWsDkM1G+ZaKDi83YImn5Ze1rMswT02/JFDQFzDn8mnJ45XPHDZ+SaKz
ZA7i5FnKd2r8e1wD8S4j/GZ1u4L7p8MENHILcqBDoURGFoKe9HQlDL4HtziWWDWR7mAj2GulB2lM
kbyGz46BCcHTR5DEX/gePcJeC0lPmycfbplG5lK3WfWwHuQqbH6pH94QvcOH0a9SkaAX8RgBiJgr
HbE6HzmWutdl59ufMXvX4cQttQr/wQ8zXCJcAiWDpYT3Z1egDtHnc9QBWxEGw1WxjtSyzrZzatA4
wCobKJllwWRe4vqLPYQJvxjYTnNPwqhh9N/fSg998tCuZ7CEpUR3TAAxosuA/u30CxNLwG/fEdnK
SeC7kflZvNLHDW6OEOSDJ8VyaQR2LgDNsbJ0UCeUas225bOt4IBM8eYQ8TvWk7voLAF0baR5X7xT
MhLZdoAEfje/T6liQf2A5L/u8pxNgE6V9HYM2Wgu2G81N983yM2K6+Ia9IM8N873bt64VvlccKp4
a0zWFrTpTPKG7L2bp5DoHf6OQ3oSJ//eZBR7CAdaVDAMj7uxI9GEaSJCgNwMT/Ad96LnXCyovur5
ZYdi781OJLjWCat+qOgF10UFRvRPoIVrS+zwi5bWhr1DeVZ/mbIq5FxZwnIcNUMG014K56f4nzrP
7u5l7332pNXGn3fkC0VfZvoZjCtltN9Ndr4FiD76S2r8ORqPyN4fcFTp+C12Kxd+0DwrxWXNxmzk
M9jthkbwr3VE5JluYJkdfXHtCcrHb7R1MYNTZZkU9kvoMBbLYDwDku6+gtJdmKimKDEW7lh4D3OQ
dzzmFOBHx7E1O9wnW7kMGA4W2+GRMuGhs3F0prZwSINgc6P+IKn02MKFH06Cj6Q0gzRc2JWgI7Kg
6f/SOYnjcDeflz/fmZ4Kzy7maKyf+FfQjbJfGkXvL2N0XseHkMqcVx/veFkwpa7IsuoQ/CuJ1+Uz
Rz+EqrArclgCKnH8XvYmNtp2v0ZcB7ttNf94RIev3R6QeT5isw2wTvVrQGLIOCVprNkgaE3G1l7P
wy6t/XHpzlZyIqOlyE0d1y3jcSL89epZxr85yztrTyLKCP++MpOImJrwO501iPfyYMYrJ+AKLPLk
IeVUrezzNpbalm5VdRdjkWalXkI5QOYmlbsZoojdHo5LYAoOPWvbg7NynXBzvNkP4VK0r5gpHaSN
/gkVbm7kGcWhA9u35FjumnTIPRIDEmCedl97eBKZbM8HEcKmNv3Ha7yU6grUoWqB0PBPSSo8U34T
jU0z9sEm8M8d/klg2NvSWxtiTTWW7mLClPM5WY9/lXqh4n07jZpsgxuR+WVo/dhHtntLV+G2AAW2
6BkX3WPBZB+XE5SKDzhpSNp5lwg2Ko7ynYUUhfWwOFWcoBN2CJTiegJqM6RRH0zZs2ONI8zj4uH7
NQuLHKdA9JjXcTv/G6aFTcK8U0eIm7FvEqN06moTjtDbliRdOHeX14bkLDMxTL2Sc9GARyksfleX
zopGS4gKwInB0qJ3RGrLWTod+CjhsbxmAqCSVsIV85Fd4lkw1MNTqygHL3kSWGJATpIViuuFC4zt
Nm0v8FOEItp1cvtqcdpBUyanEbaoaNr7YP6MsjoIaOr8FROOMMzlkuAfG3u1Q3jMMuf6pUWmH2O9
YfC38VjVtRBBHm0HPr4x7XJfmzgCXq8Ilo0tRFac/6xQHrPtT1pYVNspruyB2Mevrxcx4qkfciUn
7hOSdZmhuQWuSpRoF8VHb/kK9KnMEYolIJyFMVu+z9w+Il0kWRYuI2wpr6f6XvsTSlmvAGtoDzZY
kMQwgcsQyAoYzSp8PHPpim7DzzdNDd69NVnBwg5egPepWNkROcKXNs8PZ+wjRRYIKUJASXJY2LQR
n+asRdqfo3s902T8Zq+OVxBou8Ld2GRdITHVo3MVf5aGo8q0JkKNm3ul13FDuUoP1DfFr5RAskqu
dDfyZBWeIgOPw0v/74ZGuj2U9OWrUboGXfEZ6RWehHjmsUwFVtCh5h8uUETMgy6iwN3vJa++dymz
YdQ8RW+TlunW/mhqKSTi/JuZrEVUAsQcm3oJRME0AIqan8yxfeY6DswSCxuN9rMxD1NjLVI9ao5g
1aje7fOHC/SBLzlkIev3G8SAvFmOaC2Uz/X4sp/X3kXf0gWOjYev1BXNUa5ck5rI29a9TFja1yet
iN0fK2XL3TW80TgzHe4Xw+4jUgKIqmzOh/wvzow4UA0IEEQv3gTUCbcyNm0t1SPdo53sLfXcYQnW
DfAglAm9LhS4A1z5pODsx3omF45nyD+KvNoygxvwLfbwAvfH/t5AHekg4Ld7A3fOsFwFWLOaSSse
XCrSlQCZJKktR10N0gsHR0ohu83yujH01Fe56aytYEyBRP2QcJkgTREXNVqOYFntGFgtJqhFFTBM
k6Ncc7XMyh47DQYZbif1bMGErmvVzpV/vBifYNj4wlDM4pclbPPm3BJQGqAe0iYZpdEIBfreHLK8
CNJfwuOBYyZWqtIga+pfmPEZzSq65HrkSCPpbMc6oUe7nkT6sJVkH7ZWMowVjBtOS/xYudwOrdSb
IQwbSSvEbO99yJ8v8izSgGvGKtGv8xvW8JF0TsBKXFRiNNF3Z1G5cMDBLEb0XzZ+lCmm+NUE0TO7
M+cAe6FeD/XtG7VxXXhXzO81CHxvpKnyD4yJYReMpAw8gRk8oFwtRehCThUtfD6dRNcSy3E6Rr6I
w2Lrw7pgDeXu3EVMqk+wKWcjlv2r7OfCh9RBQhlEz6j5tmBKmjHNCMX3NpWUYxE76WoNk3+SeVIB
CsdRYZ3Pa/2RoUpJHkWRbfFxUcQMBM72ILI4QPqbnhoGo9bntJY3qIm6ecR1zwwNRedPzb9q8DYG
w0kjR3HQhLTH+lYaEDQNW2XAJ4M7jnQ1Lpl9WsZ7v+0mxIjaKyB+9RLrChbGx8jBMn7nPej//Fw1
D2mcmnEZc1G3z+x0xi6z8i31oAtF3gd91sORSIvyc2ONJRsL2H8ovyW3DW1wSQn1fJIE7BF9y0i2
IWE+I7E/OAKq21Rz82NDbFkqc0oRh5FzwceULxeaWu2dUaFQr2kX/XWxa1Gz2K/OdFBvRB4EZ1+f
F1paaLmQadnljc230cLJUoCpzcciML/sBNTYQWkv5+75DUKnjhiz86I0YITrubkc0q7f47oFW7cd
soVhYeszIAcgx2i36pS693yd8KO90LCX7FrI2HbGgh8SRRz0J9NpqsBNQME49tr8uXxRDWpOrWU/
V750cT8IjS7nDfKy4LLhf4zvLs7y84WOyZ8FPC+gkkwv34CraIOzDJ9iYtX7X4Sj88jQC+d0VTOi
Fl5mUX4wCllABtGzK29+NNODOB9rPI2Cx7zrJqld9qMpXcJ2dzocXXWyU15O0nI7+X4S42E67K9Y
Q+yIJGs/YIp+16L8pOUWtC/fgU31BiapM767CaYrXXWWIGyejvdogOjeVYz8SwhG4usZTnsPHQc5
+HLN8968ix3A/krHq/usKkf4tRYMfAPRAz3kwSXJOAZpMUo8v0QHAsx8L/NBmw8Fk9Fan1DX29ob
cREGTlzcL9lDBnCM91W8C5cPPe5m7AZP07v16BUU0U7ieYkCUuE4e3sDx6mNGajSckUnGNZqbvdK
ZUxTN0DqNKVb2QCX+6SgcZNT2e45WYLbmh7hx77MyROzzx3PK2tR9wRg1X2XGaRRFrY6wo+yI9KK
a46lliIejZJ5sN1uneT+umIIfZiMiU6XbGncqTdh48ARnFweTow+U22Wecu7VmKBNwn+evJT5Ryz
ZPFQw7DvIwrY9AkwyCcStGes8skSkEXz3cuqNPoJQNvjS01mPHyyoP7ToC322LlanXBVkZUtFxM6
kgZ/yyLLq/bL8r6Dz0ULTv1B0P8l6rcJqKiIqZCwCFwhGDzS343qrERWpMS1Y1lz4C9naj9iZ81B
H3Y89SG7KjGkUnba4/3n+q4ZHqW2tmkeTUaSIP4oxlypmn+FM0DCtskXyw5GxRkwygTdcC90ZAUa
iXVtNP08CvB7KHJcaRjRD7Pgqkx0liU2qYIK3ccyKDikrW1Ir/yvfcexiTJJ2l4Z3S3Citl5+G8f
AzSrgivZL9dO9VwAo0m8lOl10QsEoHCfy+XNVrTnzGwf5t9j6SmESV8e6GDDP8Zt6yRZUMlEZsN/
hUL+AqUoSm8lztHnIOfUP3FVLTgP1TIKv+yIX3UXp6+LTxtum0tMGWxAlayvECFnEmnoLLaEm6Yi
4AXZ0VCEq8ICrh+TFleucn7vJI7pyjRXhACiNbjtgS4jLsEPd8oKxkKAMZ1jSNuTACmflCcP1DhG
EQSWr56tkngbK4rIIrD6PyYGloae32nSFWhsSh/ehq00093KesBmHU6REnsIRqgIGi4Ul3jSdSHs
38ApH4WN4v60fUXixfq1wbNjT1Dc/f7LRlaX3pXZwJmzXCS9rmW1nK4dLm4tWfN4jN7VMFjkvRh3
LAvGXK2sQ+1E3boZJhDnti+gAFjEVK9qDJS6W/aidZCZ5q93YnGJg/R9P4TSn5+EEoNAyxpvXr3e
R27OZrof/CEtj5xo8k7FGr9yj46QigyYcdMD2jPs3d6F9yIeAShBFYQilZDUwAZLQaR9W06IctOm
4OcU1GMhiw3Du4gqvnuBiuihktOkMg74LODELduA2gmBohxu2F6fFrY+Wp1J8uzLU3Zy9gLl0Pp1
977W31SecK9GdH6qs5e/lJO3pdvpDGnA4AAfnaKGbXko2V2h0dLiwCERtVzk0xDf08xf9oYiYvaM
6SK3BXL62cPprZaI4KhRN9L5oht3a3oPd1ovmvVfTCAir1lOn/Fjr+XNMP16xQ6Tst4C/+N4L5lF
Ph+LCu//tBpLxcCRZo/IcQhqKF4eVL+YGpMjr28XHasv7ert4KypbL+Joo2WY/Lh6AnZrPHA7UHu
VP0qps10pztTMHNyniqK8EUb0muDhJPA5Fmt2LwYE/cneA3YNegB/b415g3R+XEZZ8GqYbp/T5xU
xshCRp2dBW7jGYm5CHTc4t6rxrb1kBulVQLaKrLl93OnoeCpA2vLxWcoKHXm10GzIzQqNXG2SXqc
5B6hkmhWiS+fmhV6c44WDtSXTZkakFTXpBUot+9c134VAzqmfTfADcLdpEUffkYbMvoxDuC4YtKO
6pg1Zc/TRC3IQyVSHlQGdhZ2dTiusg2CXt2zy83loWl9Eo2piLZojyX2mtZ/2ZwfrVtAOwjfg1uO
MHE/mvMKkTyv0Fnz14kjW1FgddMyih+Uhah2E2NYStX4td41iBY3t6DzwSND7z6dVXFbltJKs/1P
z+p7JEfEzZ0PTf6J448subjiaQHxQx/+5pirr2C1bByYjEk75sxpzbvpYX8HZbdqbR+gme6drIfT
J8nN02daN7OMANiI3YHPhaqpVH3kNHg+Jr8wPGERKykuATAK8uFuUtIp1a3cnYc3vN0Kh0sXD2PZ
yXBjXvhItsv35Sr4HF+zPRBDZsaq1w9Lup3OcYcJWwedhS0lsUdlxdd9PprSfG4PA+kk51QgHnPl
gWAk058A7eCneVjBQDRTbGW8QGwhDvobVuQ6GeaRSnoTUPti9CYBUddWBcRDH8z/IUD9b0jWQtfD
b477E99j+iJd0RnO87swPnoNaiVSAu49FaZo4fI1r7qjOEhlMDgY8am6UD60O9bPLNRLMF6h9IZp
1vTSJhE9Ol7OM9zjwHJtlgonZKppmT0sjzfcGPDkWild7SWRjhBb83pVLXScPmFLu+NnlCYsJhlH
ant8ywEylRXk+RAydOl74dOzw74/Eg3mPLxWyaDwjUpshYvwXOcIqvRNLjHbwVgDFMtEeK45G+bu
ir6EaXAxCmQ/vXUeIu+OWIiUHZcOE5nzlytQzQSwTWtlMomsQf7sGEqQiGhNaHt18M7kdGGXbeH6
4MK0OPhGUCBEUvRKbTADKUhaMhJWwEhCxO8srrJBibRQz9veOCSRHPjYf+dVnIM2Rf2HKPeC0nbI
ZnCJHsSSIuWtUlrB/lwQ4XkHQib9wCsJNtfduG/aV27PzAncSDV0Z3IYSUkqrN9tW0oBCsQn8jv8
vgMhEMlWa8JUfy8Pmst5Qydx3eQo4rDV7+ojGPV1gThL/avBQRoKJyz93XL6x2G5LWGVF+KsO9M0
uOHg1r+KBzqO+yjraIJCFXqxKFGWVPpCAiwQHzaZ1W+FtAzTlYw5UH9D7/G7mXjeWK4HLd+Z4cw8
9MHuVMABXDDb1W8dbtDawARXxdlJXJOpdqZUb99z6Bn/b3RkIKKh4IaECHD23ODNi0oMCqDbhuR2
U8xuGWG97V+ef8rPy7zRRwUaFlVdSjz/CLF15V6k7e2+pm5fSHXiP9jeFHIPdu6fZBpkLcXe3GpW
dGTJC/lQwT6AQJy6J0uCqt9VIH2icZ5VLFgo47PEnMBMCiA9AvrxBwmgFn2f9Kimo0R0OVuPIU6f
uqsxyaUnHoMiteMux8ENlONbm6if9PfOLRnFUrtyoKV64fjFvtLGHmz5euvB1x7bGCuCE3DTCycT
Lxy5t+7U8QY49cTOhlwZhRT8b+F07Aw+iY4cwF0lbzSb29AwnH5CG/CVHB96boyRjWkqp8aEvX49
L3gmlHz8gMFKSaKd/mmuBicz3u8iXERTQpDEH0ZuGP36+K+ZDB4UAlNSbycE/OrdFYl/XFwfTEgs
S3yiicz0FYziaPK2sV2SCAlC8rj9CmqNh8kdEODtq0YXGa5MUdStmzob/OrhbkYudoGAp2+ZkMUL
939pOl3AFKPFJKz1Ag7eHV4wXqkRZItmbVFL6tbaIM89s/PXFH4JhfF7bJY/NtcBD7HsVQMjg4DM
NZxBGb607vjza4LZdI5LxbXZ456mBve19spjJrDgYQ/mGwFiTUZLPXKwSD13LD5aoEFn/cIhdC9b
Kr3tl2Cdz4kG4q28MoNbNcijl4HaVY6kj6gt4jHPg7dn7BanjKMGKXhokgrRGXlbIjrxHQ37byh5
S/EOjybVMQSNIFTKJUAd+c5Iko2dVyIhNBuC/Pp/acdajc7jNSNcHIX0h3s4eLEO83PSJewirJm6
/nkPGgchgwfKYhPa+WmgoKLzaDhkIheq3KXMITqZvPGD+nVObwVPplv+ltz68K2BbmHXuWquJvIN
FMiw/GGC7z6VqgE/1Dp7ugbKWsgHuEwEFidCX0abhmgUvSM53g6nYNemXaKfbv85XKFqDA33hUEZ
vv4ggpSAGcqTMxWb9IsyKYPPWBw0dw9/CWVUKWnO+4/VdRzEIfxiKcIIXYegcLOo5yJZuxOLrQnc
pPK0F8udCp0FEQPpK5EVgKTLEF0DN7zvzBA/Tl9sW0+3ebw/jRbxKkCDgkH6smPKm4aPRDIL9ZRy
85VvopdhGIBWGI1WSN/xsqIz50gaya+1MQRYnPaPyRwGEZ3wtzl7nbMjsFiMcbdgyWwVIR+OkWak
M1PxdWZTLCsP+jMckDKg+MsXLapdHAWQ9/PaUcWsMBKxEsXvLwrfuxg8QhpXgJrByYwN8HGnG3rw
V7bzpj0MQg6pxGSDzAbLqXHESTHKC2WFKQ5wxXMS2BGuk9CBM6T/HtwoeHRG9gvEtTQnzpQgYT3R
hJbeyGg/E91uPkdOHbOq+OD22UE0wJuzHtBgwD7lq77VqDNetBsheZCyUy6BlwJkib41k4iQ7/I6
POo+Ylq1hHByMDTc/1Kzj3+90EA4SAgWFQLf9blN0Pgjvka8kwH9qdT6AmiHxGOrcuEjwklQQmj8
Ns9fqWMxJU8XrAI4sdUXpls/wCEnEAm80+NHNUMjQNA0WFVpw38qHPYK8OL3nG46R9Jr4Z5WL6K0
oYVymNhJOBX1LW0Exd559HN1hHaprtNoYAlHz+p9SpyOXUEwsqUyX0xlFiSzpj5fYcVbDDMce3r/
QoNNIYZXpiTlaPF0wFJtOA/POTzbK9X8dKy9hC3QMJRU/UaIjWP6htgi0mjIfvEVOfT3xduBEKCw
iK1Qf2AyaP1w2XObYYf1F7jh0TOMRdrak7u+BS5ytGb/rpqz/4Rlnaou1cM0+12DHa9yRFPiEsAr
9VO6iu9hY7692i+wsIPQBXrJu/5AxY8ywXcRXlCde1DWhgfUZ5dd0JlCQDcHBhznpOx7Fx6GTs0v
LC/54HXssXME4dY+nDkMGFGUaKs75MLOGDIGvatiLFmReDa71lpgKEhsPGDMZBKoOPPkCT6mIwKx
B7ZUIAqsPdNdyKm7VSxmksfOqW5fTkZeq0/HBSeUvLDY2gCn8Vef6FJV112LyI8yNY7JerK+cri6
uEwIPwudHEhBqQ9SPvrkNbGdCz0n2zCLsSWcSa5tcf+9enp9U7AZUWioM5DbjZcHlt0cG3vu2c80
tNrA44z+69asAd1nR0f/YE3yr27D01UOb34HtP3n3l30a/4x0qdjrX/7SH16gXOzqAA9VMiqSogR
6AWW7iyOf/w2+12UXLQoGyC3p1gZgyJONBiE1BI+x9VKUYsN6Q3MuChoklgKznOLG+Lz3uSCMYNy
uV8bi39defiUE32j9jTYIxRgM4X745XeyTyU2VEUWvP3MOZwrlGpTyeY9U1pDjSX41W3xpyRztKM
TkpV+UKF39bFnbKq+mhpb1Bl/nmjoNznRpiIK4ek4Z9OtR2dX8nOcvJt51sIU2HfLKTUP/7lXXJ4
mCGgWRDcSij44V7He2b6yM8PKHmxXO0M125Uhw+XiMiPUqXO0pGCusXU/3d8CzYmSZtYGXxwKWzM
qgXXw1wJR9w49FhfkNGF7Uz07M65UgOWHtkGqX0O/eKww66kAWwSMpPmDT6Yk9KEIeUXWwv8pW8M
kFaqiJ5Fo8XMIm4C+7kOyABdfIFGVfe4+U7re/RYi6sv0vbaCqejG84a3xZHuEM/8CsiVyXk+/WC
pEKNE7PHS3BPfRWqdapvuYM8aVGWFzb9vVhpEb7aDg2KmkqoY+tnv0MXk3uJKrMtyK+oywmHOJwN
IyNJs/J+HksprQuTrItxUZyO+WA57WNCdCJVJgnEIcPmMPrgiAoI5RQ8lcoSCpRcLrCE09nLMyQx
1JFI80/M+sXJV8KeGqfQBfgi+x/XBTFrmnkmEu7RlUeOShmRxuMMhLAmrSQ2uwVPp/l4aXu28FXN
qWFjCshBCYR1rEFYquvNFO7lSkzQKIYiZ5WOLg2M++D55uQUJVb9tRdP5nmnvQekzAN8wOJMPUZ5
RemGlkdXMe9ZRBq/FV3WrFjrGVqfx5seJNBtDIHFsClLl6VO9yL+4gVjdAcSRaZGa17HJHV1IJhY
SHijv8ABf/ynyUJ/Ds2O45GB16E8jt6JxsDkOP3GL73YmAaG971Bs2TcK16kL7n+VAJDmOfBUorT
D7x1vbP/8njC04p1HBuqP+/6ENvZB88+v3XxNXLzzDVQN0X4OjnNhpcu8MzLuqqvr+1wgq+xe1hR
+TIpIMtfl4IzNUIrfs/qZzWiM6wcvQFVXZdvgOsaE8BPkHE9VnHM3qs5M033mvytkZBmth0Qooz1
9G/hHOYbtADjo9yPo3+R4HFY7laAtfZ9DffGGoukBzN47H3MzAPepzJ3lWJBw+JZkTtCXEVWTD9b
1NgJ7wFP6Y6DxGTC8wi2qaeTldFJj+dXB8NCUV98aQ5xz3i1LSPiU1cRwfc/86igKNicHSTseSrK
6JyVoHm71ED+IWX/YrP3e2KB+xHyjEvC2a9zdINbTsJ8cNb9cianstZJz3960vatxWqwoeSV+8oL
2lNZge40HSJIFCk2Kn/LdcN4lPQhuLna6pQCtSCQej9jtJfK3mjhAmZ9gdxVSja7G0r53mfocRD1
jqYFyZAHXVrk1h34G5Sn3OCvEM0doIHxyrXZQuwMHnuvdwPVrVtG8LzbnPMKoyoKRYBnLc1w9bP9
zuodpx3Yomi2QA/SGolm5wQ1sNfcWVYXaDxCCp0IGT5uT6lZboML/5nctfcI0p6TRH6SstfzqrKc
H2ZKev0PWaYOt2nRWmL6qODRVXiMkFRw757k3BYRoVh3nm8lJ1ns+1tmmlFJOIeQoj3jt2/5nP2M
pOx5M7mVBCnVI5o1XhhdJWB4LsuAc6FSuT3JSRtZoyMvA8KFpd2in6DuNqOyfj5BJSutSS0PpM62
AeaqSaUoCTEv8sn0kKDxQ2OHZE3Uuwgk1xwdn1xFYm2A32EMIC13pwYcacAh4IM13c1L5R4tDM1Y
8VPANOWNB6jlwgQkjxKRLlBoNk5wof24/gM0ewyngoX6E3cyYXbwKO4wK7UQ+6NnSgif02DHiYWa
5CCVoiHNxIGhz8TBGXkOJVIWiSxruR5y+M+2K+0y9ZDbLMPF4DgtpCBUE1HcVZWxm//ctahUp3U3
ZfRpMJPFKJn+GGESgK+vEJtDV5aCcnRRqVQmxkX3kRhza7mgFA62ctueJrz1NLcZsazxxrg8XlZd
EnkuWt4z6UOKDzCbtl8wplAOeYq7Y+EoYPYyK/+OBuvI+h4l8sP8IzuOmM/6l6VE8BP45XETCUKC
edWpwL2J/+7lhYo4Lc6h1w2KSXEiAmWX0gWCG8bJ6dHSaeLqsCoopXMNfQmWHETp5J1qz5a0NaAg
29HvudBs+pa6EMNyU4VvGhhsqMnr4dHOItVS41msbfH13eygMpOx314JTIm5hY7IQsgGAdxvyFuF
q0T6AXujaVlzgbeD59jv/hFaAX/rdcNtgYWA7gCc4IcUy83e0hajtvhdZW/wmIyYcuLheRhjX2+b
8E+YCVadlUAk3VEpa8XKP5g6zkSAUuJfsVaxy6HpsTJNOXgjHJZy58EvY75+k1nrjgTHqO+szIRv
tye+M15Z6ys4G+MMok7KunL24GUeDYtgdVB2IxR1aZyKTm33Ryu3+ePOYazRHurI4/iYeXYSS0JN
0MGD4CMNHdADpxOS+LZlFgrWhkrYPA/f7J920+AzZa8UyYylXOrrX3TFEeR1mK7efzEHUkPMq/h9
mrj0X/Df0AUtsAdqLIHUlFQKbRAuSkR5z4aNMuzvpVRqRJKj6tDSgjT6M/j+H3XalzeZuO2rPI3K
6M4LOWRNtiwSkdfDO1ILLAhptNP3R+VF3wwSCJz3NORa8uqw4zWwnMdWsKc8GucXYJFQHB5f9Hd+
k8+FC94lzgobwQEzkGgu2osDwnTC34K6IaZaJUVfxF5XNKa+KjemttFGC/wPKqYdwv6+c4/lviTD
V2Tok3Q+mBWC9cHP9Cl+rQ63v589mn4bgFEUjuMEzefUi6BJjE+xOdYWPOGcBhDxOLsUq+IHuNtA
C14XVFPY2b+RZGFpNZHmw6kX9t59pC1zQrJgvtkg1VDFshOoBwa+ED2sBUDFxdMu3V0HyTMCV1y8
WlprJwCzQcZZ8S3WQj4WjN/lpV9trwzVzlhK/wNjXJvNTY9W86uoaEs0JVdVVEWgE5c+RHJA2NAY
Rq0+dqdM3lqIfCyXA2/p+uJbBj4oPML1rtW9rkFuEO30izOQT1/xwAP1lyEJcTTfsoWVgiiIo0Ao
r/qz2fSTfBmR1cY4rUJw6FgZcayBgSNHA0051nSoEyJhlfP79lAuJzUNPwI7XBNawNioBxPC2zVR
TAjktepvkPvV+aUgJwVBehS15rt5XHc05kWLYq9Hd2hM9SZpOwaKWT2xhgx0pkCB0+kjJDvmQbQi
0qV8D2QIWFmE7dr7RG73cHoAxttQ0i1AQsY/BqDofbM6Arrt03nfClHHy5zj9mfAfmIkTaF3EFKF
TNzVTswrcsrGrHcYqA2gUq3nnRZ/9nf0w0CzTSXx2GQYwmi8xnSpsfo7izZ3KV20xu9CWYigcDeN
QksQBR4cBinankcPhefxxW1Ja4fRezvkfyqCbDxUt1rwZQV81n120D4CZCa2fkUSGG9d/9c5niY7
KcAc1F1/RGBGTXk2iqhxGWplJ2KyGhpzeoyx+Ay/Ks//18l4Z438/5LVF7T53X61chT2Vulnr9SI
Sdnxal1HzVnpo9V0aKWrLBjT3rg+FkFx4AP9FnSPLb5jAUT46tGpf20ojxzarpFn9G3H/azjA5Dd
4GmfrjRFDRQvp3wWlnqkK3HGpMMKhbFrrFzM4UTd/85lKF5n0eTQtN7g2Lt8g5BYd0qFGrYl+Xqb
zpAFOrcnuyP3zOCZUHvDiVIcACXI6qKTS53kDPc7btMkwCXoYAImmitxFSPJeD8vYokkBkM0upOj
5iYQH9ST8H6PyPbg1OXweSH9HruCgXwXRf6HCQua6FCyP8fCowozfwGm9ZKJM52sf4lYaYT6/TiC
62XXyLnCf66bwgmszy7vMpMZurawc1HXuySE3sfw4OQH1nnSLEZBweEZEwwI5RBo8m9DT1rzLeXr
Esv/wEqkYKt1mnR2JqAhzmaVZWyJSPnYIyqoRNVioKBpf9RurZzfaGYB25d4Mekh6gOQx3QvFRiG
QmhHvdFnJHTaLMDP90Kjh5B2McX1WVSngrXlUEET9jjea4hZiuqj2PlXL+Mnp8ajjJSu+i3Wh9lf
D5bDj1ZwoajIC6AF0CiL9PvQQka28DVlgNMzpGmBnvQgHr5Yjadn8wLlKBj8N0lYSNozggPe/Dau
GLpw2vB3ztC9WpW25YSI2mKXplnDHOQGnmodR+vNibOFOJnC/RdJN+kkWRU6jOY+1YUqDHXZAPoK
tD30EHXW25GG/z2rY1XaY+edPSpc+IzlPPUyZpyuAfGapWMnZ89FweIDj8bjQGbaohFzNv7kTaqy
/jKIivWKlyN/3BWrPM9nzz+2ma08FRxHIWAnWe6ulUN7s3UcBejBOY4GFCODYX3ZvXsQmnZp4yVe
Qw8Y1itPyD0vUJOlhHHTteMfXRUByMsHh8DKV91uxUmCsnn7i/zwAd8PWUTG9t/QgYAg+gFoZ1/M
QRV/5ZRgBgr0w9Bv4d/qir9VulJmbXKpFXDc/adXi10GqIS/xWUqAY+c4Cq00HkefBoQDOG/xPrm
CLP344UDy7Sw7CkFufwrztMynS/oiLPxoulhDn3dcOUq0UqJuqE/CGCHBH/cLDdsYm0r2QCcympA
wbRMNxZpNsrXKjhtaRKjQejJKYt+J4WpumBlK6t2xRYqr2Zw7KZDh9YAbyUqYGC15/lpZjI5RRij
bUlEX0iUrmz8SAAL29jLqvtCO4HxrQU37nXHQqq0ri7qst4S3segXTHRqVFkNqSgmznRZ+dL+kDs
GY2xipWXVtBqxjaw/lBR9EW8JmHzPk4RrxyX7TC++E80G/x4uGem15BpM3FdzK8a77rewbAKR9O+
zSkweSnGxOc2B3ab0tRlcZVQFMF05RP2Ht7PVXAFHdpl7tHasF6uS0CV6uIWvIt6qcpppnp7IPvL
NBnwLGMxBw6EtDGb4xPn9jF7L9DPpZx+vG43g+At6gV4Jjxbn83X4I4C4WPp3MddRBh4M9AkdLzX
3+mNujAp2CuqfKCPB8MgZblXJquVv1Rxvi1wfGFL7zCdM9vrAUo5kwGTrbD1qxxRBnlKuuxukhxy
xv2SRs9LY2whk0w9xiFUKUgOx3Bl6VvQgYsBUGDyzQ1EkYsxrbFyZIihQpKiOHzR9Z5ql1dvCgiD
96217ji6TrHi5MU5F1bnYaEMk4AQA6JMBaFkjdUmYdh0ZKr6LvddRooQHNqztA5CIDuM60FzQj8x
NfKk4YxFxKeBJUKN3v5lTG6hMal4wU+Db/AhkAloNLqZzVTd2ruD9ZVIxb++DmZW10Kpj527xAaS
/sjJ+SQ3YgyxJtKpeeBHzU7bW7x+xkhtP2eDpwSjt5fYUAab7FJ2tcuVesd+6NSuc7m1KKfqrEaD
GnZ9yXzUKff0IJG8zZW9lC207KN0i52NFRic86P+tuP9kI074iix+KgeGBTSfaLcojlu67N2czFa
9Co7K2ffbw6C0+UGEUOcSeiGfXBnZTRCJKYhsW2P3WCVr/VRFxA9xmKWG7yR2+ml1kRW+YgNcVrL
uMF/WUBOlgjVgEuHNXbcrSEzbOuyy/0/C8aeMFVad+e7FrHheVxg1/iM7XKsjao5R28XvZVRll9P
auAD8Z77BsTxhLSW4n8dk6FkKNA7DGW1mA5SUGqTBbV66VkpgedSvj6aeK9sAptfaEO96lpwNeJo
IxX5bFF6iWTs/LIlMOg0E1xk8UwXx1xB73N2dndLFLaRpuGWTUCSiu697EH1/+dMXxu6AQZYNik9
Ri6do0xp03NVKKZBmem1eEtGKG0pnWGpeMcc/v0YOOyr0QHNJqmw4ahzv5xzNOfAN96srkwmUMeJ
QalTe7gt51bO6ujVAHaO3O01nXbaHRu5pYKFOqdRsSD20B2nArc+tMTuCCtrhSwm7JwqtUo0SrZg
YmIigz2/rSmZ0fpgwa67lDUf5gK8QdN9sMU3aYR2HfYutgml4JztRuBWW80l/ZFQHmMB5bpWW9NJ
mh+f80l+TmaGgH03uuupjhUVOjM/sPCIWumvwjQbT2YT2W3myaqnFMMbytFuvXmi9wcLRwtCLU7d
DE0f1/obLhUJq3NhUjX4Nio78AekzhBUVL1T4C8vFugY7p+CF0LtOlhB9F1UzUteGAiub+cktHu9
japV+P+94HdIXFe+5fsWDyoGd8nsYSmNsMEakZ039MlrNMX4BRqly4LUAds9Y+hvWyMjFWk+hRxy
6tGcyGm8HrjWG7h5LB8So1qE+I7V3utGWPbRAVAX4oszGNpzAYSeXovJ5rYCCB5X9b0LayR4Gjtu
Kn/L0PLSJZGIkdm2vil7TnXB4X0QHN/mneCaDJpf/ifr6AsRJVelsHzULzPuB6NUp9vjHDLTJT9q
rY7+Lr5I1AfYkWUzfYfX+aYqCBfgHt1Csy5/SrYUU7ZhKiXi3Ag7emKrhepec0lNpvyrOn/AmGoh
DtmSgRv6eCHr4Qa9OMNnWey4UPNaWHBj4/xe8Knp+qaUvEExVOMfdU8aW5kD9W9IoTdc5udAx6jY
pKk6OM2HdfxaqOPrX0oP0y8S2XLtgQsYsb+Nk+g8MTtXdT8cNU1E5Ti9HzGX6zHW38cUQvW7PFYE
2+lM6xU6+lpgHEDuHK9/miUENOsbpK4ZtLw9gyLqq+KqdlFDXnOykjTyFDZiuFMcQ8SUU8vFQxV3
SEvcBZgUDn6lSqhXZbGiz2dZWvjb3Oa88UuFzxwCUXcP142j2KELxhuRAwokD4oVAxNHRhhUApjY
iiwszrVEraOcI0/Lq5y+0sbzryZtxxGn5JwuEGjbYddOV7DpY08O9nfyv0Szzz2xFsiTSZYCyEQ1
Bc8DExdk9zGzWJEXgsbhlozbxTTE5FJJEewkGkJhrHYLHfd8+/8bSoCascCtUC1uz7bjDIxN/gkM
ozPCU0jEId91gN2oves7DK7vaMuAwGvzdIPGM5MQS8r2lKXTGF7TiGQ2vZ6nG+VmjlWaULSKBjMq
pKknZfOTFNkgrGvM/jLh/TljmNTY+yP+8qq5NfuXkC15bqXg3FAKV1lF81TcTNdjE6A1IvHqN0WA
AeteQKDdPXG47D2wcE70gVrHeFBs7CGC7BJQbBayG88w9kOw6XVWUl/0fnifSZdpgjqOffe+EkYZ
1WZ0EwR2hTlhhVsiLYD1Xc9gXuywMb38Zw3R6XcwsH5yzGlAPpJHPM5qzNtb9VvnSNIPyZ2kqgrj
9xm7eLQvUmLGvAdDniFYno4ozvI92C3ambKi9Lfk1e0kd/3WTAVowfxPJTX2Enopke+hf7K9ou5J
4EFrsLB0o5XSiY0nasyGjvV0MjmNkFX2MKIZArPUaBqUL0hPsiIN3s0h9+HGuALA/iJRz9htlgWZ
l+jbTDga659qrwLopkuT36TaVx5+LWxRPRC+j/ld3C2qU9wjAosjj+5RPqehzy85p6tl0/igZrVy
qwkL+68Rnfxi0Qw2zTQaOTSPo2o3PfW2FjRqN9Gef2O4IIh9HG43z2Ikg/jI/fKRSJEfUwFrhoU0
pFPy0a2LIYQgKPEhQM/5eu8AFAPddfWY52ZqOArIXL3LY/mLxgVOgA7igN9PoB5Fb8HTOqeJJVEt
dkoejT2cjYdsBVdpQBSGd8vGy15f27fqYtuNwp0Pb0xA6vsIDYfpA64qgH2LGusBEWUaDawl3lZr
zaKdvZjtiZzVo72PX0e1H+l2cKCjAqd60WVsx8to+Vn3N+FeFkiYSzqVaj6sUvsitoQuwoGI5pBr
K3NS1nTyxrU2zX0NlTny/zPQ5Lljjjj+f16LElKgg8OIUD04RvbkIe2f736km8TLPWlcE4mERVwe
4RyUyB33Upws1F3Et90VTrQDfb3p8DmRDj3kIfYZBRZiD5uuuj3ms40N3acqbRvr5Qxl088ROU3A
JUwRu/Jb28WKK7mVn5iFJoW6LOtQn2usxm4QgS9MOJ+0xnxugoLA1AP4Znjey5pLdXBOm16+3R3/
Nx6Hb+coFMEE0S/yIveslPuiz9lAoYpHIienHGtFNhU+m8CNt1Mi3H3lyZVbz0I0mikgswcnDz+n
ZCWMdU56Z/h1BaBtZwycYnvZ+d9tAWY6F6jjx154xxmvfPRpu/8BqjD3fJT1a1LTaZugTBXe7c81
vskAfo3mKlz+Wy4xb0RMyVt53XRfACYWP3MUorxJvCrz8ULrxqka5LxGV85fitey6AgwzA5rFDsB
B93nMP+OY89SybvPNPrjktbqe8lo5Rngu3R1XIQZV0OjtLHR3FjobxTw1tPhFEelFtr80gB46FNV
8U+BzmyHAEwPr0+BH5xyVi+y8JsOmrg0XZrhmLP/xMQLHPTh3Ns8BjXU2Mt5osYbFgYZen/GlNKf
sv+faN2QqPox7LajsMrJYidswcyuDpJWiEd7Jx6VAS0idclyUFjoCL6H3mFmftmHRjiQfQczncYS
qNdeADAj0UuYjumjFYx8ZdbmEbgl2j25V3FYNJgUPCMeRIEhEAKPeIJd13MNSN0t0Jg8dB456F7z
4in7IJCBmLA/ubl82zTGyMX440lsw3m4uJNDI4pHAIX3OCXsKbyt4X557D3W8oC9qMRRopIVrLmR
YkUmGMIgNlkUzlzjQzdTvPnb5uoG1M7cq3DvnVu4ANgfZpDcEMMTSeSvKCI3bQ3OzjKEWgVuYCtp
JSJRoTkVwyu6x5mQs0pMh+bSWTiB6K87jTZw2q4ncTvpvPYeeJ/i4IT9w/GrAbz6DJJW1u1wFVDv
G7K1oXtMlWaoa09AL95b/siNmBMExhCoYt9s2D2xVSAVg8g3cJrlFbmjFV4TzTnHh5MIaBpAPGVZ
lMT3LYv3V5BCGVDTjgFbVBQuoeYEakbtX9FAYOLDI8JpF9KiEsY64KXDhtcnog3Pb3qEelEYezjQ
6zMmgoPat8E2wIhhqaaWbDqv6D2mY37fQuTIHDDBsE6UKfrR2ESRYBWVGCGgXpt/XW09W2VjPv2Q
l0ze/vQe/uOY29OF/cgmgCR5r92KwVSQ2ObLAX8hMBl5V1T70Y4KfoEj4WKYBis2nL+2EEfbBtQI
02gsI45qGLxmGYlzrwZXGjKj33i4/SY1WIQ1qV688Akgnr1f430AWWogjz5z7i3fY9Z1MOkK0E1I
nSzJPDI5GMytjodYsf/JHCbpWD++OrfDcQ5lN4oOgO96PalSGYwQAsjwGOzw/bQpetU2B6FcLibr
3XEqLGACAigrNbnm7d9yAtEvK3NpSWCRCyrdCUNErqZRcqZT24O9jZ5nTA29Q63EftF2M0sL+0Ue
u6h8yYe2M93b+QK0HsGdZp1KxIsStfj8zYbIPhbcPW/vZpP8IUKzo2bC19OPIKPk6n6rVIrs8H98
yGmneL5Q6hWu1KDwN65CItO7xUgPdzcXz+pOeqgwM+iHdLMDHX3EsCOmrxrc9zxognR4X7r7gtJK
Ac8KwcR33HmL2K86x8dyXmw+/70huszlbXbQdcBhLjPG9JZf70i22Ow16in5fhH15KDhcsumhNG+
AAeZ56xcv8efBA8E6euioi2JbE7cVw2ui07XAM5C2P2mzvcVIaK+qMv3tEgGq8fZ7HSoPpvo9Qx2
eD4IsxLLjkAfQkWGt+t3W0ITEM+EEFeSiDmgKPO2OCP5owEXf793Hsrl/j/X5qn/s4d5Z301Hzed
7z2L+eCxoGhCHvO+g3Axc0O3diYgi+j5xjRmUgxKiL1yRlbmecTOoRWT1Mm+uvF7JDm1Fr0k/znZ
2NFYr6fwJ6IQT+SeZ4Qjk2z8QgPnZT7aWvBRcQ76IgKz7RkPOTtVuA9/rGH08+qXlyEoOuSZk6nj
PMmUTqbEozNMg8OAtMF8UvNqkMZIQ8LEf9KOLVw9VcX9bmPlOPVH4l8Y+Oy1wBEWc1e/SApSnwJ2
ETZjqKesKDC+iwvBaZOYAQ25X1OzuO2Eckjb3Ls/FUDawSiN9VhbDTNwbyuNBDZwLxhMGsOaWw8O
Pvdk3Pt8zDflwvM6udgY2JT2gIil1ndUqIUeSW/W5fjabtMzc+cZp/vf8GobtMlbEq1AMtDGCB+i
A5+1DSRF+sK37ub8kTOQLgPsKxstpaUNfpgRCItpv1O1iQH+M0gFR0qqr8sXFzQWJJAbNm0YQASe
3FntQkCn3MSV0/N7LQRed0OOPwy5eykQHx+mDkYsv8CKyLGXUMSa2voKpGfJv+Viw2XELvRMq/pC
xzeHn4su7bHhNgKtGqSS8B3AAcPaenFJ12tvcx5KAUv81xbRRjO+NaQ9oXEE0PxE6uN8oLBekBql
oiiazEJDx2SXyOQKcVZBLQUkYyvmSW5/3T+bExz5A+vP5c5034nLEfllP2hCOMSZ9pi5N4FiBs1C
PNizTn+h6/wmYR3Le9teIXRbjwqTzog/Gmqcz6GUZFTLFx8lUomTlZS8S5vDeL9ycrHQVJM1K/3F
NprIHtLVhtpe/MtqjFupl99cvjdABnYP5489c6SBsclDV3pBBztexHnX2gyKFOfYsV6lmc8/fkPP
7c0DAFkF9FNw60Ozo+Mpo3s56Lx76pfVBPwdFJVA/N0XYOPBHTHtEkyADevKZzLQS8GpgNkweIKs
BtsxGBuv8sJmw7faOaTolNSIMtROprIGOxmZRPtrlzTZN24ooTFmp5ahISvYjiVGWqj5k7FCQbvq
plJKg+iqAce/m5mIaZ8W/t3wuHl8oQFmfQFRCSCwi0UlJrFD4PjohnphroYtFXdLwi8FTw2I8Rz5
HQIhKuKRQd+pI1w/kHYrfEdNDs5PnZvt6YBN3lhs+mFGy5drdyuS56silZZAVMHPkE82xSSUH/ge
6C4aPWbEZBfxYriEo8V7Eo0fPKxfYD617b2UvGrGGfnciNXFcGxpWTriziJr2LlHZGLGGIrskuob
eBG4MO1D92xRZk1XmkhWrD6R8PUg7O8nE00qpZ85KpqnFVaikc0e542Q2k8JFUvmY4I81DpY6c7v
32KF/N8zALSRZYWZs1L8plzftLAKoDUpe4xDfVjmn+e8YgteITdvl46ia7sxac3wZRkJsOX6CVnI
iX0gM0zl+KpsA1N5xVGs9siJOQlpX8+s0VTJT/iq755Xt6z0MWqJAgslAAIAIUPSdspNwIQE8FAQ
E+XUX4pkkE8LsKQUA2rCCk2N7r86jO5UrE5WhuKKkySaWamstSjeV7xq9UxDk0wRtKl4JLGqK6Jg
Gjh1uzX3Fs6EEkuM6vtenWysWirC7B4f+2IHolZgbv62Mi7bSeYFjTQVC+Kz2wcNTigqG1+rEnu1
8+Drdt2v2XRso3ZHRftQYp/d6wA+sU3XNAiW8AziIVGtjLjJPC+Jad1SAn9aRBPi3Q7X3BQ62ROW
u4+KntDUcK6sAX6qd+a6zJ0HBbbo/7g7JejE+gQHLiLdtDWCMv2inBMbQDmRgi9L30IhRTpA15/o
wFOq+Q12DrUHXGWLErLhmuvCuiHlmpvF6oI29g9EL6JSedOWJe7EhWz4/g8pxT+Mi7ukg4AMjd94
yhFPRDVHiZe46ymLJTJpdLuAkm90VgLrdJDDS4cxnoi3JbWxdti4lFeJEYxPJLKmY1gjSzDZKVTO
ZaKErP6zweLrcR+cWym7brKzMzj62APP/6+9f9AmvehR3sMlzksSoz22eOqWyxyt5dsxBlc6Ih8w
IpVxT93Cy7CS3uT0s6ZGxFnTxVhUNs1qekNEBuawIEpXMYsl9pQUB1dxsGGk6N45y+duOOVvVAzs
+CHvpKdWFBfw0TxeXHrVVH018jQhrN2D9pBhSbnvEpsz8GOIzmRFOaGgt8w6wDWwi+nK2hz5KIb1
HEMkB4nW9l3PGOLW7ZhbB8X8MLHy0Gdw44XaS5j1iREUV1EBeJBWaLHiWoQHYJnLWsoMQYW8txz+
BpKI4xWW2efyB0RlTkv5+4EDVtsb4Kq/g90szeDOmkV3mvihdffvk7ab9uQgv2qq6CnWJQODlMXE
xlZwRdca5GSpSfSFqgHfw7AHKfzbwdJyeIEK/pV9ts+RDOvJHeC5L3XUeegOF+S3CWWCgrmSSXsH
RAQrRk9YxSVZyktWDosjjiyBsH68fMei3/vokGyYSaWtqiNfqoEvRGt8llhKVVeDXIHkZ0BGF8JY
rip6Jq1uM0y7EMN/S2VofkoNcqgTHM4BA+JIpNrG59ZKMBFEkXUpVg9GnR4bsQZV+8ID55gqgtJC
UGpm/BXmo1hv8goQxLwk9K73p0r1M7Ukzf0TYBzlj+lmkHDQuMeygiRvghRVchU/ptgYoxogA8K0
GDnysYz15TKQZRXPTaL6RFV6aGg9rqTbjtpIX8tgmMDNFJgFgj4CzSNUf/qkGoS5eshzCdd8GEj1
8siC80jMIZ0Tq3ktUOK+e6MWeMi7wz5/3vEFYyz7s80jHwj68Y4UBpe491gzYw+5pkvSyfJBm2aZ
ucM80ww0FZJpEXFNXMfVtkxRCtqzPZJo5BVoV4x3TnvNqW6/BXaJQ5b+QoEkxKdB0w0svQ8nQjgc
i0t52Wssp/soT6QKYr89evxA1wMjWT+pEZ/nuPYqJtrkThggqSrEg1O1+tLsuDNzxQugBHy2gjZ9
C3+zFeC9Gq8HnTmHFlQ9UqOO9qPHKnrFwlWYe/msN9TCU0vsZ05vMldXz9Qr03U/d8c+C3EUv5q7
6s3K2A1jvvdE4HeOWl5IFimhnNtxBGYFQ7nkWd1lgqeIIcM8q14dRPYaVBgqG8gZQYPu8b6kw0CH
9u4eFNuuF5FUbDN+p7hwZMsTif67hjvyer0c+HgM9h5bnb78Fo4etCoXs3IqB7gbexTbvYaXDhWd
xJyMtTVm80qnT6mTEM2WnqgWKpmuFrwr4K0d792ZKJirAKHRp13jiVtjWH3U3n8OtztZ1ULxmYVw
cRVVTl0/OY7HT3APEZJsOlYS5xWWUOSDoGRGieBpLLjjREPwB49MXVPA1f8UKOXAr8UhQzbn7X4Z
HAf98YpE5n9A4PtAGpGqxhdjRSVBnNfgEfNdiouC9DzRVn4qyK2jfbIGJhiiKx5bPWLhcAl+Jadz
z9XdteuJfDabdsZfdkk3myHB7L4FNi9xr5Z4I8gIKfAbrmqBAcW9GERWfeUiuhi0TP5u4MbUkhAc
4Z1xyPuJNkB+OqTc7uOOm2eECUS1IYuK6vEIx9Lq/USF1V7ISQFaunPNSGxUdPp7d6tUx905C6cP
pBRT/sZhD85f/2KNhj6KxOxL5aZAXnqNtdvwctUubHbHcEBlAOFeJ+kGRzOBZBdPG8pDKSCZ5qql
89fjrq/b84TJH/Qa2jheDXxaJ7hhWv5Tv21/mRkbkiMd6/uyhtabjtICb7z+orSxelEn/kXQmZoE
kqwlrF7rXnOwECs4s55wrnGxcrvJ7JVArswBChbAnf2VgjubL4ayGVCKA35sm8yx6YGb0MG8Gr7/
XIgkvW53Ia1ZUzFiGPIQShutUYC893PY1+VGjebDk8/SGBEHXnVuOWsBJZgbWBUdbTHGctwYNTOJ
ueVMCc8enuj5iXmsgjznK89MYg2fptBsLfWgysPYvc1iXQhumItmbq+qmBY76lfeaRiZE2eAlsTN
8iscvQUC2JqFiC8EL3riV0J91BHZe/ZgSH0VSsi8OB8ePjJ1oXUYI6ZwiDkw2aYUcYvSfwYyAGmD
csx3e/SGoKM2aBGiVkfGDH5pIhQ0Mxf6+kGfiq2SZcMo6wvJUjTSfxlVdzr28ffTHNHDMCxCnJMn
6Hcwoplcf3OA1wr9P1schhu1HE5yC1D7kovQ0IFnwum14P52NHC70c1XG962WyDSa/jQAq8zPt2i
MKw0UZ4dc8hnkujORTPZT305wSdRdjVnyaBUODUz/2fXK9pdKNwDTKqbCe0DDs3Kvey20cJwePZ9
nmTAFWqQXcpF7bN+meTfw3EC9KVh1sYbEDPVN3jlSERQSeVtJ8TyrdHkj5LAHG9ZO3Jry6ARRfLm
PZDcEYtroXD3+RJZHm7pfn0oD6S5SYBqUYxliFL/mWFHRzXQZIj3THuhbOFnuUpGUakzcXoLOx72
dpfRAwoMcbktOPPWAvWmmQVETeiM8PSiqeUKrhB3Sd+y4ZZM/DFSCq12KnoDVi9yHnhp/SreveIV
B6iE48rxPHOoQTX+hf0UUz+ktLp5SpnRHq2mVvOH42mL6rzK+x17FhkNhn7PhTxjCmup9G/+ksRW
y7KzFfqm/NbloopzmVFt4bQa6TdRbQRCggBR4+sdVhSHA75+Gh0yq6J1qrfYnwzdz2uSmw23Ju6c
OTYUm81qP6DzQXeX+0S+G3WDJAAQng4V9nBRURxi95tt9VAkUYDJmnjSdADxwS5lczLTg681Jhqs
gmbqgW+2vNzShCgteB8ODw9aQgLlhA+she0peY16iazK+bgd+PgcbO+og28ZZ4+GhSJs6yBGMAqH
Rl3TXUZt1dULz65hMxueU2nE6xYjjNkF985gIFTK9fLQ2Cp1PpabZCleUBKtKZR0kLmP+wZBM2US
heg96BGyj9EDnajMsbvYw6IGz/as2cw1i45oO0aoepvLmNNGE5mbA/dO0zEdNXRt1QL57+0Dum5y
cG5q5bd0hzml4MtKYpCkc4SPrSdktBEx79b001e9gUePzM5lYIOU0WR047hcVeyOJEUe0eBwNzmY
9tAM0ymfMp7DakuYKjC7pqXET55ktdDS9SgGx4jEYfrs3YqPJcbNQg/faYd2sGWeLGDutjugTZu4
mms6MLb030alDNlhuDqhIMWYbyGxHW/QQ6tvU4gKCe8By+OLVXsd/uWSx6xBqOZyIuF6qnIex8fl
My1BoduFI9DvHB9zjV8APeujEdRl6+CbdpCz0xSRqvR77nY2OuktwwuHU6UFZtOVlxzXJN7UgBOd
G/mXsKLyUl2aUB7xuMfyPrujusr0IYZxx+k662YOg2V/KSvf4g83M74gCaoTduNVlzzKi5hHmqcC
/6LP/XAAhyq28/+5aPsEvVjCMuR2hIOi3lD0OyXT0oKK3knWKrsonMnT0VqH0IpXmGmdGvl44wHI
csM8ajmJxpyxCvDaUVQv0z7K47kPftcOkxjxPzmIFDny9TfyQMqTrqFGVzOM67VoKlUTvRk/M0o1
uBtkq6vDYtNx31AOitap3md/yRpYuMm09ro7gaMuG9uYSC64QhXL1u1t5xe2ye6M+lDgSenUDlih
S3C2b/P0SQU9044NnKptGhtWcF7G91IKHAArbP6FUpg/RfmIT1ZS/54oEdqecEwLSZYGiavTyNiz
t5GMhymvVDZ1okWbGcX089Eg6PpTAw+Q9lY0/Pt3+afUroQsPs8FN6/LSWjSpAZtyrzPw3Uqwp0D
E+sp3xqFl3rdFtrAfI9LLrhlA2AegrsyyYfqhNgRndUEzcVwnOEPbNAWMY0QjeMxBUz40iWfZaJA
dKS6UWuEg3EqYcHSPGaoIoJY02NqXCkEsyL85DbMA7Lz5zmsWW0QYA6vXrhi5Dh5Jw9SWHHxZW5Y
GwEY5TQF4ULJ3Q/JxkeNmgSr+wYWRGw4tz/ZKEDkUVIYhxL3FYQrHDwo4gc9QoRKOk7hQwxcplSZ
MePB0+GwD+sEraz/V8hUSvm4pdHmdeslNnZegWK4jP3YHpH2Ss0DedfTX/HeFJy2UhisH+oa/HuX
+PLCwwqTVxS5Z5aBcufziqyj7hbDA8Vc/YA+1hlMD+HizdmK1ixN4wiNuRtx6EVHQzdT3KkVQgfS
rmuRa5HoYHXVEFXqicZyPaqFxMlz/d1KDBm45Z8RJlZiAmsyBQYavBTikzaHsEvlP7TqgvcSjhUY
vquOzo54Tzb2QQvpJkqtHzCh2ipI+PHk8lNVMxhUKSTm8744jHmxFgX9SDHnXjzkpmbpwLRhYtGN
n94qAQzpeF44KUCR/E4Q4n18DhfMyDKhosiGjuW97tdA34YvoziHZBfqlp3S0/+SL9p7gPe3JrBm
x9ylUG9ZXa21HkTMS/Eg/2Z7ANCiXBF/ERHcsuCaC5AdDHi3uGqy6kuK9O8F95aA0YMgucSO5xvs
hV/hpXxu95FbrYxU8IUmjBlLnadkyE0n4OsKlHMjtrz6VBQ1YjurZGkBePX60YJ6AnHrXobPVdwW
OzSSHDdlU+b7azyL4Auwnq1RbXS4B9W85p1iWngZd3rPkD7m0AC20UQxgnrFqChpR2ut4wfWX9YX
K9hzpwtHaFAI996u3Iqo92+SgS2ST7hivJuyUua/fRZDDS2QnPcxV0MxDH0G+EAMaM7K2m90PYVk
kozhNbtfMnNPTy6YfGtXYLuRTyuLmn/d7FeLnL1JOCFGHHJg9C5uhkKHTkHnlD8k/5YaR4IlGrj0
nfvhGeQAzX5lFE3d3zU0VO1JiSH2w6yJT0sPIQzzV4AI8ARkUsLsvruWuxP8Md+jKsyZQJFR/EZ4
OykKbw1xwXEtORBdVLA8ZQ+uqCIeOPoGarM2diUB22C0P+fqPNgo3GY+sypSG9HvqOt5iImjRPdT
1qr4sExLX1EJz+E+8O6JM0u8dsq4kNprsSgYDBMBtUzwBF5JoETjIRJqUXbauImdEf1SpL2xbpFV
EaA/QpkUXpEUdvoqfEKxJTBhME6gc7yaLvwyUVxbSUobOQuuGXW7OBhrHb4GnsLMHA2tn7L1aFRQ
w8voS/XdYWbAPbJqYPblWcSHCOGvjPjWcb9QWNGZd7/pvkGTEJW2lk2acDG9gjsjLGdr3p/TLAnH
IXLsz5V2OKtRlwO+J3v2RFkycU0f27E06eaX15c4362eCP+gbGy6/xbFrXhgstUYVI4aOtoBfQvb
0nRmsvA2j2TDwr6Hij1WbwGWS/gLtodbUJXZfxVUw8qjTZjCIx4JOHkJjhAX4kN6wPjj+GOSoJo/
vYxn6LuuRrZp9SM9entflIGa2y11yVkUo/Gzt+3JcCjrJcOLjm+l+M4nLttErm/DB9IvdOojGKpp
WB/GVwevhLGiaIOS6HkDQdoZxRD4GisV4k6FUhve+1XaykmAs03bj4JsKEmQ5REiOodnnKqZsoXd
h+j1LZ/I7I+icSpvOWQbadd/o7jjDClXrymfl4eudayF97oFnxHb/4rTDt4sYcrp6hg8S+VJaRkV
AfMskM6bvGWSLpU3eHHwB8Nb5IzZzkRzQmWbWBrmxWhofq125K5VUn8rrvHVxKY1wmSrEUqqfByy
UXRvkxdl0kb0tAjfpMB61z2LZpQUDg21boQRckeKh6O0AbpKXrgACsn9oxeN4ydv+URiQn0l6Itc
IcVvo7m7SDszLT9vNfhQkMxHJcnagrqfpD/5tP74HONJEEFjvDhBN1gEGbsAEmWrJ37TYCyTinDk
8I+FhV02ztsfJHPuZNRJGv3cQVG+MwR7J1/AFLQE760R9XuIGKb/yvEKoqwP088nn4opiHjX3StP
SVOIzK4wKqt9kvmwiwhH6rvjgO5i3gIXGS+yCXOR1CUSo250gEEbapEhwcqMtW75mWcJBSxmbHpu
QGepStMyGTWn+Y4C8eiKwiltThwiBhCWZ3FHWdU2V4zxKWwlAcoErPtVF5yEEzJX4AolPnmin8Jn
bSNeGS9VhqkTMC67B+VaZCIN6HlAB3CntSawhFkYDL6CIOLMMQfrzVllfDqPk0PzCCaOKfCGxSzp
x6V4vCfb+xdlSDZiF/fV9r7xDRmXElmkd90EXUgPnRi6YfROughA2iqqzWOu/GOSQe3Z1BDDpdfH
tLRX+JSI2MoDJCjdcNpSluJsvUNZF3A/tLg1GrYQ8YUmqPzbUSPo+XMuVye+wxaSpdcsiOmsYQ5W
f3/YaAGepp2vTE/3xNlXHeiSCUoVsR44kLCdDx9dVTMspOK1dLa5kbCT2sKloSvoaYkDGykUIK6l
+gjCS1zKtEnkCofsCWc6AaD1nlZhZjLLyKc+a/p/Wbww/jxKfumXntS27Gqihp+/ADZ5DJcdt8/E
fAX9tJdcBmhm5EcM5k3ZZJQahBo0AfX+dBt2eR5CYFhugJMbC0ZO4fhl7Kg3TNyxsOBJcecJpWb2
NS6sDquRbmCvriPSC5k7Wquiz5CWs9shSnaAJy1hI7hIy2QfPPYBj+YayslTwAJWDEAcsXT2wHS9
1kD+MeJRkDBorvc1R76ijf2YVuvuooczLcvnMYFEdpfpQ0Bt4yYAXA4fS3pY9TzSCJgD7v0FOryp
lmtTZIN6vMnQtBiXz+SId79oCpPslhOEoDEFPJR5ZEcZ6RBHAaiyGKER3ASCsCIa+kQt3z7L6GVl
V+n/RZaLcoNBkm69RnQ7Ep4ppDoWwRT03ufKkFwiOqot1fYvBaIc3B5k1WWWKzqNRMPGcLkX4WBW
7LWq0B2f2EuqX/UmZgnHXYdvOev4nAD8VxmGW/3X/1HMqKY3HxFWNvqVj+Vtk0I7HCTAjqgIxjln
agzYyHKqVKTBr47LEW6JswI88lwQ3KMF0HVqsPhZwWmKD6olvpNsP235o4i3iBtkEDEXYq/8zV9X
fgYYiE9LwSm5pUJU9UmM+nACQOlHm7xup+hvo6HFN5TnD/uX1QqWqmyS5SpZ7m4hso9kWKQO/TqI
PugMubLR2VKouPMxayHVDM3V3TLr8Q/+9I2HTvBOon+4VZnRhCgJWraPtplB0+7iQS60GVDZWOka
QmumUIXEgGtfeEnwrW3ow7H653GHDXnqOYssmRzKm+BDY8SR4emhxPJkQ5zAxAjnMxLKjlbzKT4f
sMJsjZA+lTFBOuz79gC9dZJko58Td2qOGaXUp/4fJQy+qcQbxFlKP4pq8DKi0JkT1Yw+hV6w8VDJ
YUYyMG/mVTYsuDDeuMa994463dPsWJOMdFnudaLuku/dWb0+gdhYnqGrvSU6AoaztPOwEWjpeitK
uAg1L0+tI/YEDqOMpLWZYi52XjpQm4JXlpD53+k+0SLOoSZjiFpiksKO2kO8R5w7dmUM/RWxKXFi
Z+kh1/WxfJNN0y81XFcwDfEUSkqo36Vpp8TdvkZYmNT+aEMRNZjDRT3ffZ65oGKPk3bJmpFMy6H9
zi6Y5cX3QY9xzuI2IkroRP17LlaiwBno/URjSQgulplKUlENf4B4ipU1DOhprA/1fGvNe0HooJNi
I29XdLl4X7eFMRchzYMMDzR9zcaKDPhLSMrnV4vI0sGRa6e96zKm0eeTwhDK9otDTVaS38KeDU6C
pH7PeCq55rxfe4nvAtdOmneBDrpM1zfhBaANYcuxQWmHaO1TVLRO4/m7DVquw131WS0URgHGA+RP
Eb1IbEVcueQFX7/vQkPSj7bvyTE3O1xw93x1bBC1mRJBh4EQJ11drcaT3VCGFBVfDXjETV/VG3Mp
xNOS3cesaa90QPTZlIYAbzHE5vCs+GTwXnKPnEbB6LdupdofeqUAw6EjNmUi1zIm80h6F+UpaSX/
v5P2ZaW+6dUq1EshRTrAJsJIsrekPLLdi17wT6NaSnWd+6W+d69oCb68CUxZdk86mfg2SE/n4lCP
Ty0XzZFjHSvnqlaoa/kQOJW/ECnhln0D8YcsogMwhswJbZPtGpwEBGMmL5/x0CEEv2oMwAHCnr1j
bvvnlQsl/eL0K5GNRiM2V26rUkYAuoAy15BIJlbx0slodYax4Lp0Nh1zSv3jR75T2/3pb1jNhhKT
CJ+01ap5td5yUmuERp3qCjRIj5OYavIK9FHl1A8GsHY+UP4CRpn5qK0+xhwwU1FtSUF1dukMjVGA
Npfp9uvvYwF4PXNyTzzvqtzWNQxDEwmu66nuCswW4dXg4JpKXSStjzYbR3Et7M6LNgwne4j74+iX
6+YygIwSRXGLSNCptHO2hS66Mtn4AJzahx2FI6769aCkyo1GyoXHTqEhV9uoNqbEHky6axzzz86p
KOATpcvU3+NOp2QBFlPf6d4/WxyCnM6/jq7Irp3ZEWyz81zJbDyNUvXGfFo/S39aJOlCin/CxC0b
7mQ1i35LI6eutj5B/OM52GUEmRvn707EsO3FU2/g+KtYUSDKcdp9XAF1Akq1gLG00iJIS0LHAVxk
GvjOMTcYI3EBeEiokbiYADzHIW0UWWGtKdVKom/oqadEtr+y9XkmGMjMrQVUFjKH2yTHn1legpYg
WVL12Aoqr3HEqr0z0wDX13n9pcMAQqdka2HmkvckdKqAPxKbp2raVnKkTNkbhE5uwC4ZaqKyMw7u
f4bW0hkPjf/r0M/G7ZmuEI+sYRoGIb6FlEFxxdIs52r1Pp7DS55WwXH/94/A81W1HcM4Or7hhPQh
e7FbksfFsw6z8hHP+eSZ2TaPLZEkQmET4hxQV7Y9Lgb6BeACQ8IecXM1fSh/UkQv7W64iEF0arA8
3lYcp9vPkFOxcN09vGF8HE2as727UO3coBM7zVomZGZtgcsyl43olxuzWZOU4YfHYrC6cFOrlZwv
OAZb9eWTrXvPl5O50o3BhSTq6+vYGRxoHMvgcXqUX01dJPuvT1uiUhaY2bxOKW8+27Kd7tUjuWbP
5uT13ZZXM0XnYMkHzQlbA4ygw613CQ1LyEo0JcOSr2QRA1Nr7drEvYvtarQIC2CQuaE/spiLNWBw
ZdNP4wtZGRBoFpLkLgPuybjhWkEfJuqHlaRqvAVfZGg6zDfs40Y4zbKLHo7A4B2216fJvrt+ImcD
z+T49xHrncT8HHuqfEe1XSHUVx32oFvhs+fALeb3Oj/3XkuKxFqgd2XW8TR44rsbKbkDda19544H
wYJV+h8CD9V4B20PAP7cSv+eY34K9IIv1Ozoy9y5B7U4T5YnKv5VjmNpLrcJynv1C/F7+XazJn1i
I0cO/CVFa7fj5goIPC+lB8gfqxlKbiyhcf+cKaPMw/HMfcDPQupMHPPTXhLamA/88i7XkvKnVEd6
L5Vb5RRWs8tbwpEr5byJsbI32cisihOlfSqGhotnK81REkR7vluMie/bZYvKEe+mdKSEprkBqI9O
PwmhVRWC9i4CvlThr9lFl5f8E4Kxmv5SMCZpxRtUcAhqKLVn60iY3sTnc9Ae/TEdLq8XPUwWh3U0
ffLXE1ej4vftBXDYXmMUt/uYUzA8tGGNvQs7hR5dwUEQ4D4IN4zvw3oYdXW3tNFE+9E16jJgb3qd
+QYqPzckO7ecektjhk1xPGZAHKUOqssN/shUZXyHKXXPoarFMJDCZREIpOaRQapIAQFR0ro/NYVg
UxStjlGclkbBDi9ld7EEMYyVNdFk++/0OspYJ/zP6byS9ArSm1m0CWCzm1Toiol6FMswOCT4V80S
j7VUOL8nXPtIqTFpxn9pACqk78WsMx5CNDn0Dx05pplMMsThlFE6shAQ+pDA9EcfPUInwFfD0/Qq
+CP6FuA//xuBR5HsqKmaO2sP6/EU7ZM2OmS8NYoGVpXFB4QtVBto3jKFIr4YVDadz/OHpoWYpDaU
pys1U0zoqkg7USj1McpLBUq+xCocUDkbzJUIei0Kgk6cg7axKoCmoJthyRvjkD3/LKfTNzjG5kjA
l5WjYBmd0rgpmC8zgq90xzQ1lT0QF7k/AjBruUiqiAFkX3thYJ5OpC/htIDj3XpkIZ8vyhGjxrv+
qoU6hFvr7IWPHutkHIF23f6jD33rrjk++KbI2jGbtcvNHuijYxw5NbdawO+xkTemVCjBkipXbnxK
2aHtNkhowAiY9zsjiEispLrauSt8lzENfZ6c+jpXfCMng0qsll5ula5celb98FfI4Uu5kwUjqtTp
WfmeE9Y4fko9zp4WK5J9LbNbV4TPLEZezJeuYtz29A0LJyHfMRfNxAJIdoYLJWWyPKcllN5rWOt+
S4CBrRuvwF3Nl19j2aLVwS91dvv6Fbb1oU68Uh8Z6k+W9l6OBN5QsAxVMmMt9OlvAD8WMrIMT/F7
zYXcTUxeUFBQEvNxTiSf8oQYGkdau2qrcXp1XX8c7z195+hScRO7IWI48uZvM3mr89m+QVATGYUe
Vj/+RsiJnvSpqKfjQZt3lxisRWnMMnkECLcsZxZKi5dnoSuerCsK3sXws7jY+LDU/rpaGrE97t1d
RFy96Du/AzTx/dVtuLjI71InriA5cw+CdcNpk+o5W4sRbt/VBVMCq0WLhC5QiCViviKQtjmD4Wa2
mkyN6S7KFfLzK7d8sEDssJCZyywA/IYe8QpJ5U5SI+wtjtJ/LyMtQu+/tZFSNo8mQK9jpo1Yq+Iy
+bkrLbkA2FfRUYb/LGN3Si940TThtWiItLBZMtmDxH4b80YZgTqD3xhlS8hcKgGG1DNsHORq9Unh
TFx2eX4Ro494mlnsTBXEdHblxRjf5PBEpVkaYx8fcLFe4uQwQ2MZ8w3gudObarz9Ebm8KqRWK8R2
bcssuk0c9DtXt06BwpAo+rhyuJ2QfZ55PYbEI+6s2UEeUkVZLQUJulSf+gV3Llnm8t4EBwhAGmXV
XwHfxyvzcvraPriIiql1pqmjCDGjO/nJ3j2vFZ64jL6iEdcLRo+4TjnDf5/zb1ZThaPl2ia0nk47
qx4JnX9QpEat/sfVP/Xbh3MQW9YFS3HoGJG2IGGwVhh0yA9VGS4zkuU+R3tl4YPHTVzhKQg2/yy5
wqjl7Hl+fxnXQzPK1Nh/Gmj0/vbGDSHjDkBdIaFdq3L4fHsrI/9edus1oPnTwsm/EuzJKfnWb+SC
HDhBD0jEYQUoZ+Yc07MFxbGhrYUZJ0s4P3YwxvIhdnPwxvuk1AJXH8FKRB+oR4iFj48kJfUqBGfI
zGvfR3i8+3nD2DDMCk+bQcH4L3u/SRi+CGV01LzDS/RTYlLShnGidsq2ARFblrSQJlDtmx/DhqPY
WmjrQmFM1UiEfpIVG6X2bjWI+a1RN1mYjOcujHlEkfoCp+9obaxpvY8mhkAM3hXhtba8rC6gghoJ
CieP4Mu3CZDqQkQY3g1v76J+nY2l96p6vUAjpFCqNF9Q4VuwySZJxTyCCLehSjcYY10vk0KPBfAd
R5T5P7k8azsongwzH0Xn9AiciCPglwu4z1BPym/blJq7gXzldcFukPjTpM1RXlMbPHesm7d7Y0mi
BtPyIaVF+5ESISu0qQ7C6ho920hhOs9dh3qQum8M1LvWw9Cd2Z3KMRdogmDuNHesaSHYcgrepZlr
nEXrMPrPMjnid5CjBxj9ghFSDjq6CI17aotY7y0WWSFPrv3F3y+C8Z1N2CFORarJwduA0OVUDCQ8
Iw0Ni26U1PbBmzNrRSpPC8A/z8Wq6UoXbyY1vScQTH1Kw0CTXoOq+MEEosHJb4wrwVk+u5hEYZhK
A4mzwRe9GbHR+EnlarSQypvenNmAg7tmo2pIiJoCTo98mD8kRuDPiEs0RS4I7CUTke0x/rbG0HZI
4IF47HtqjmUpT36c8nAjnG1vohz2pnlDijvo1yB+FaUE4LIrTx2OFhqHb7rAo16Nld9DZ52J60xK
zoCVjEjZz4Da60AehyMc8ZA4SfN+tMO3m18FILk2kuS//YyRdJUnhFTt7J+uI8s5oGWtqIlSqL4J
G39ZUkrzQPnFf5e1TdvF8RiJRQ5UvFPjj0y/dE6uLEgzdR52E4XUKuD3HsOIB+P2KHH9wuAgCblB
yQZ+1weWoBzBks5GTc+l/Ws0cqc01Okvkyp03h9+2M4Oqlf3Hrp93r4J1snziCpguDM0Qo1SNkQh
Mces+JGoFtH0YcMu+kmmjZ9dTPFA6hs8bjTI8W3N+0TEmEfcbmBJfezaBej7IsV/QQvJee8tz6my
FuiyI7hf9VLeDNMKKqTfOVmQVGLExWciaPG3btdZK30z2yz+/pvjrNqmaghWnDDH1CYpfZJe+eM4
yM7erWFUumL8ryM3EVDBewHIt2OEiTZ70kECorkp4c/RzfYMXs7nELIe+Y6essKrX+8tKD+inTWh
/UOA1zEd9Isd4O9PEFuv3hzrfE8uW7r91YmIru1/xo6q958vuyb6fpnmZEurE2dcSoBhF1icZUhI
8o9uQ/JwMFDNd68oPDIazgp7eUZLp6PTRqOx4DsItJrew5+yJQ2D1G3UWnNYO6xHRzJlml3FZVZF
WvtlokMYCk4g+avhwHRjsUdCOFJJCAhO5fOcCuwLO2f52P1DLOmKtlGknBkUQ+4LFqo7RkWzRYcA
u6YklxqRXz42jkbvlkb1wZkttHIXGlT6Ou7FdlgVOcSsx6hVoqNexPgn1i0xvor2C0Vm+6W6a15U
I2Zg4N83+z7rGrlemll79JeYSbq4ip5loj4wfs+qFOZeksxe+9CYmHyizPu2GlEQTvdhSSYF8ZVK
EDoVPg8DJFrC9ka2Ao6XsnQHxIhxxlVA9PNZvgHswryZBZxfiXEXqGOPbb4RavoqeCuqKpBafTI4
1xxBjE9qpMZp069ICCaao+R7WPH+HNTTdW3F5L2LdDLjIV/vLSqxZhFWKrQOeCv3kV2Y+S3TEg7l
DVZogURmsQEYWg8ut8Rgdf1aPAJsgjpI9/BNMffb1XBUoAx4vj+ZifYPG+Q1TTUCgTRdkI7aQuOs
5PUDCJ/1Cifunh4xohYnz8Wu6v9L3nmPlFl7ezj0HWA5NRhw0n5pDDs5YEqoID6GM0iPmb0Ps363
Qqf8vUdVzsCeX4Fcvpeqz8dqD1KfssuPck+0Y0fOv1tJMuRBfw6IpWQiKUwNhungPdC44FqjoJ53
N0jSRndFG9g0UvhtB3S/fBGnVm84++ZKyCvIbqtIBuc4i2pVxyixdEPo1aszxveZVcSteuLvxpxl
4DxKvzMwp2lmShl8SP+5/VEEyFgw3Fo+kWKUgGc65ZI1N1mVJn6djGsy8tsQUtamSYBLUrnndjfS
VSvKYzHfyNhVKRmrC3mrDauJbswgwBZnToGVrIXReCHgs9TTb7zGtvjGP80YX2eWNBvYAK9FFpcF
VCo+GrCiXSiDgEk32oYmL4pewVwJjlKRiqEwWsslaYdBXmsUnkI4VXm6xADxp01OONB3nDpZpBkc
Fcb+SXXmgp9qKHdUDrzU61APAo0cGf49LbxDd4wU66je2/BeBwjVRtYI4Eqcd6a2IuGPWjTkRUIK
ZlFNI5ZI1AmmOjIM8dqAyiB6pcpYD8NDrj6b/Ni0qb3bWq4Fj7rOquovfvRhXWGAFgAiHDfucX2u
KXrugO/Guqu6HYnpeeiETSDGGJHKFqDisoY85k7WC/E7W4D5HVyd+qSYbSYO04IdpeZGQ/ynP75g
EFtzpz3kQ8bbJ4dzNPgykF/ND1qPUIuSyRoHeSW+nrSgX2OdznHidoCxaO3z0WZwPNwaFP0ywA1i
os9W9aln/V7va0qKRPBBXi2BNWy0qbpj1TJmUBDuGdEq73w3QVvWpKNTmAVfJ6yOZltSqFS6szE4
R9n2j+RY8EaJkQk9jFHvuS+xrTd4GlVfiNfyUi6lonrXxV4omb9kSoHrAtMI8mUXe/zt6PWPwvmf
V4zj54TnkYbk8ryGjaMmlW0F1ciZnPxRiI0i+lTPh1Ml1ptNF5nvEIqUFe4frjKBBhZs3DIRxf0t
uZ5Kg0WeUKte3zuxwRYPC6ogLGZif5DA8kAKCh/BxsvLzWwqtBJY2lAEEUS2TXLpvClCkkjxZuGc
JTuWGGatHZA6VhdQ1wxXAuBSNkOLGr1zTWHil8b0sVVcfyXicXLycJaMqs+i6Rnms+xJnPFlznv8
uO06S/nwI1tdxMflFRSlPjXT9q9ubJsUoX30M+gkrS1cYqPBe/VUz0rcu3JnbQ+8iq47q5rd+Ure
2HGzJ/HebD/eku2TgASuvr3Z6XJ4DQIpgdeHPCicQP0HNGmj9Mxjq+QRD+qHKtBneKKBQTtvHDNq
NS7WhV1Da0PUz7WKoGn34yj8g1R4vK6hh03FGKEfl4/fTskpFJbFg1S0FO1podVCZv2GXCS6XovX
V4HEUIIYrzGVWhtSbSIO32kFv9Y5WnIK87w2OQruF5u196nLg9TKlCP+eOSZGnKWvom8Zej0BH2Z
HPAx9R16egCLyGkL0N6dlYVQcMX3zXUu+548/QuyPad+O5zau4e3eklVczuw2pNpBa6eJrKSxnkG
CkqU16UdrMXjKIQGPxCxCCK/eka0T8USXyQ3grAvj38ziONM9Pam0T8Uz2m1nJc3UrNBFJ9CZ5tH
lC7bIEEOQWPcPY1caa+0TfF8nfhEV1gyN2DpENNOk/jcHnVnxTPv7md0+Bc9wYwrk+GDCl6X0dWI
QmWf/ktRoQSe7kYWJWqyExo7ETxaPM0jLZgTUoIrtr5Pjn6z1uTFCxeu4QXt65nF7yQv+vgtKEhn
I4+27e8Mq3wvO5spGWUw8GQXdsxVkV/e249uPmWkwg/baqNvjLafRj8fWXolG3hkNBpfxjjBQ62X
v498Bc7lKuwBnje8OIvHkHdi3rV9/f+2Ra9bS9ZEtf16u+XYx3cpMgqZyQbQAvnVbRg7wvBRS89Q
HtHS7cW90wp4alePa+JTKb2khIYhu06eyEcHCj80Xaqy6ywaHYXvqzXcPtiMXcSrTXoVt09PcOO7
CsSRsZ/J1mdI7YS1WPd2MC+X15KladH9oA2WKdDzgbuSsYwnfYV6VWetbAQ26FJGXwv5fjUGJyvk
LUjLyYlMZnyon3ttzm6offbqz7+uCISKh/T84+8tm+gvKpeWXfGMnjJwgdfXYD7ZEbDLzj8xZgLO
xTEh/KDgYQfUZDP7kUdlbsmGRcfpLFU4xgA+ipKZIHda1nZoFCX7IJ8kkgY0/7dlDB+g+BWVoEEi
C822TIXVDSKtXwU0r3HT/VabZdo+swHK8PyhThwlNrV4RbjswYRfZkDqfY4NF9Gqav6Cpkc4iJa0
9tRydGqYsLemqGXmiKWI0OnNEK/tMJO7JY6HuMvTpYhESWrpiFP+zMosoTaRtFRNsk1P/umVDIOl
wtVXMyEA3jXGHWlbaVrIwTlZK62TxVU7yAMkC//SXQVTWhIJMJxqw8zkuDNZwbY9DzlinOeI8sVK
GnjclZFuZbRVZew0G/BjCxvQvif+x/friW8MEVV5bh8kyVyUa97RX3NKlOG1ojtw3UOe9KyXl3JI
bs/reaR8LjmiN0kankpoNOhl01LjDQr75rp4wI6S2FQ7SfBWYVtBgIv9blP81Itsg36AqCrPVgsJ
fefMQXQ/Zx1HRWuyDXAkYkJKk4aimvPD6SkBe3XoN9KEjf9ei5PEvjkL1wsAbWhJn5L/A4Fs66Ou
MqnssKQVb41knXtOJUQH/5ZdUB18A7SvpMa0ZufbwsdE3Bf/Aq2bNCbrA7C+yjg3g1lUhTp9YMre
/0lidnO8GgsR9am3BGhBclgHBPZFyI3TSZxilvQqTOoFPDaT6OOEcqs0FsfISGVg4fHtoogSosIb
q8fkzl2kYuFkeaTF+sqg3YGUCEE/oOKPxDOLc+SVWu0SIeMwj8amE93vOliA5oMtExGyvaMRtV7y
kP0A8AL6ykxewk3rI0ntDvGEaUPvsrihw/3Qiw4O0WPKnQ6VlQi/CihBRi/tHh5t5ZMUhAqwC/mo
C45tCSTndqK2zJDHWQOIOrZMJuvXEO9P9J2deQCTh/uzwMOpDZfkPV8+Nixhh0jJHufGxvG+r8NP
xYQdgQ5/C834CBZkiu9+MYnG5kdv7Z2F0/+eGe3nx+YhJmWMJHBa/azixEBN7NlGGuG1wtHT9AdH
Tdx6zO9hV/E/u4ZWrdzHQFo2m9pVjmCNa0p4ceqA3CwbNo3HMLpUkxUfyV3FzDYpIOqn/fqNHYlB
oksrLbzI5pMr6fmULx+21eQjpeS5Uo+BOeYwsvzhWo19Q2UskfRinWONH9xeL2lIZ+OtM6Oy1FgR
Ua4MpKxo2eUCPAvUS1HlqOZ5ytBgU1MuRWY26fHOlOUFaunoNXwEWj3FsWT5mNGoTLa68gW8ZrXu
wCZFXsB/07/7X3htq8ncc/UNgmTVCi50FB5UMETjqJXUoBEGBqId2KvF1zC2gd+9DRs8vyMlpa/v
zXdqI89W79suJabMPlvPchLecSqBojpgeKhJ3DrnYF1qj7XnFAZ2OGfSsV4Srf60EyByCMhyOqXQ
++DTYYCf2BtWGZnXGajnuRQebIKtUjmHIPoR3n/Aqv2Ek3u+iDsahrE8e3RvF767m0aIHHDOj82K
Nv4IbWCBwnUo/Vkuk45yP78kSExU8RSckuZxooH0FmsnSWLDrpCYhQgaFAg3KZKb3ou9q323bc6p
0wc5jCrKvrl7RTVsfJPnggF+5H9obiZ+I6+59DDyF0i3gU+yqq3gE+XdAqIBZES1s0jYGszDMWfn
ooX01L3aeFmAYZJTSEMdxtItl12P95CdAtYED2z+tmVBTSMiy84QWINhFkwwFVIhqbvnZPlxrsL8
4ZTz4kbZDnIrAikPrZhnFbI758TBevsYqZamZ+gRlPxa8sxQOI3nN4X6Akv261FJOCdCgb+Nm0Ok
d4dCxPtnh981tB5PbMtIqb8YGCij0RuJZwsWZfJoqCM90rHKRk2ms/ybi5eP/gm4TsNTOUCh7Yc4
gGyt+4k84cFrZXneRK3lye7kUMzACTpJzsVGh/rCt1/a4qI4fzIzDL7Dselreci4ulJjXSzxdhzC
nzeIw8XvFicYA2Z4K2RoaZsFcgBsSftxhIMI+1useDnD+UxGN+qjsGLNLww/SwljEqgqEe6fRPAZ
ajcUuRxred9OJfzgeFNO85pXx38dQuZzwwaRm2MWsOWEfuCoGhPp6uk85eO+O18A5aAGW3SbRd1S
J3TbWyvJl4AxCERjnb3F8KM/g/dYByMSmOMXT5gFqZJ56KhS3EGSwDiiLpHpM9InX0APiy2Dx5EJ
gDdBs6y8xKsRqxI5ulOzIdE6AtddvEjUS6ENZnXLceLUobQHQYvqXaRiotLTMo0EDVIpQzAy2t11
aMcHaKbNksyteLC9oLpOQ876wwr9CSg6GAKtBXJc8EUgH4u/D6X7biH1tSFQsiQFhtMqUPrFWcC4
QTDeTCN/7jobEX0gIIR+OBcUNadzlKwo03UOLUZL/2czdOozLPHvehVv8PE1UHRzZ2S99uulghy8
fLKK+V1GWVMhwHMvPoTLcIMyOMJBy10N2qx/no4yXIJwYsLA3E/nfwTDJn9B5XlmnjALmn+P55gi
LIwIHxwyU3ki0FKNJ+fxnwfP+pFCnYKO893fxdyQbp36EwVexMcysFFtjnkNZlltteS7ok/7t5gu
/hAoEjosJVqA8NtNc3GAdzFR9JNgPcTFpPiTPlleKU/UM1O9i9r7wokFXjI12e1VPN+qtBytIF5c
0A32cJgl25gQ254c6l6yRNVFvbOp3wR1YXQA2qsIdjXjkcTu5BPqc7kUimt60YTP6qJq3RL4h3Gl
lDOpzfozNGvPXbV04u1m+VcVAD8DqbGO2rpH0tk5Nu8RIQqqCbpWGJR40INxOjKovG0PwvawfEnk
LYW7R6DML3DHX264v3qbhn09XDEIuiVlzBQSam4MF51tM1ljQVJ9oGXQT3Da1o5VcHUVTFJWu7nE
YA/amtrIkSFPEzpyasO91oXtro6tPkJ/tHkyEOhdYktmxTDt+xlbjHQ6nHtpA4d5m+aysAVSmEqD
s/WHfwLUAdMwOqiaKm7ferhsSejyju9ZKYosAjer9qgMALs3ILO3rO21ZjCmEqWKILJZWBTXaoQG
fpQCnNRLACySLt01CfoNS+LoACDJTjpjAwJ0J2DANvdj+eqRAOKQqZb1A9XAQdpzlu4e0RR8bM8V
3/T5a6pkpVXd8/FEj6jfEuRnwfwFK9fJ6LxmyIk/MWJAiqRcCXvo0zoTLoh0izipnQ9o6/P01eNV
L6+qDyTN7Z4l7Pkz/HLeyBBihU/1qOoKRhg334KraALfQG3Ns9oJfaLWljd9FGRWwNBbcFesf+Gj
2onP8bz32AcHZeCoCmCxwIgv6gQokdF10ZfXSxdbnqCsWW1vec9KGL7yEAiEnOFnbWfVTs54mRs9
i3O4i1iSuH+KLfIVB8l7tQHITT817hM3ehpAc8O0wLN5ms6xEvfeqStM7GkAPHftC6B/rPWmiTQe
AwMgWcmh82khz50NQpu6GQuaTfA3cA3Rp7b7w2BYIzwNllDQL5Pw96cH/3QMGVDfSShtk/VuQifm
NFLdJHwyjq94eT3coUkB5Dsf9HIr5alqQxAom4yyxONNh0zqbNXotk8ohUuzO+93X+sLlZf9WN/S
lJ0lVr9P3Gn+f56g8NCpgQsbotUDMOeN5NBWwzWrCWz7H97/QwvTfSzQlmnlhvUorEDwqNRt2E1k
Y3mT3L6ac0X7/fgo6IDKtS7n23QHSMyaqwihytIppXieBY1Z+DXZR2Z1O182zo8dtueHqpmLOigA
no0d4aQx0hZl9kQ/SD/MC+oRuSFu438bzcU7OdZo2oGxOrkCNDfTT4wAWc6HoqSmV7gNUw23XUs7
WbGdbSVc1xkChSoHtqfs/iupr8+xBr/uKD3WqYsTvyR038hGbGXb2mX6JueZxPmt7ujNQZqZgFN3
yRozrJQtR61v2Pv/EnpCcsuYbe5enVRTWwopxyDTBS7izUO7PwuZ07wrZXQJE078By3VJT4pn4qo
fUwR1NT77ZtrTWOK0gtDA61ziggW4RkjXdoR0Ldt3c6r9rPi5tfJ+OVaKJF52sjCnBTLo8TEWG0o
1An3IKoMMcbzDyOrYMO0t5r8mcWoy4FVbP8mgelEMDNDLrx+ZMr+XTbYq/8R/lcyjFWndoAyGa7x
hu8ETUHrWKlga5uzJFosblpm7AiMr8jcnns8iNfsQcjXvodK7sLclO0XMVpJfGLYXxDSudlLOI5p
6pvCA1umX3R89ALe68h0xk9ycco0m4F2DpKrPQxh/D8NthW1+iQEJE4HbTo/SWHH6jBHL28rLcg7
Q9DZjbLbUrklnQSgRx6d5d2FCQEH0a9mInZPzG2De78tPosx0TFXLNA6yp5qMP2At3AbCMdbvKOo
Q2M9T+2Q9rUnIUgwxeCGwJf9JVQIcfEn0zWz4lKb9fpUmWEhbFTkkAiPuUVEdlZCaXfgbqaFWCS7
ozNvK3CIlAqU9/ExgHgP64B0p+HWhDlwcgR/0WeTg3aSIYi6NgMB2XezoAHdYIpKJo0G03gQNbAf
9chb+M657dK+4noK+YqtFJ/WS101+iCBynZkb+zD
`protect end_protected
